LIBRARY  IEEE; 
USE  IEEE.STD_LOGIC_1164.ALL; 
USE  IEEE.STD_LOGIC_ARITH.ALL; 
USE  IEEE.STD_LOGIC_UNSIGNED.ALL;
 
ENTITY color_rom_vhd  IS 
	PORT( 
	    i_M_US          : IN STD_LOGIC; -- atas
	    i_K_US          : IN STD_LOGIC; -- bawah
	    i_H_US          : IN STD_LOGIC; -- kanan
	    i_M_BT          : IN STD_LOGIC; -- kiri
	    i_K_BT          : IN STD_LOGIC; -- MULAI/RESET
	    i_H_BT          : IN STD_LOGIC; -- waktu
	    i_pixel_column  : IN STD_LOGIC_VECTOR( 9 DOWNTO 0 );
	    i_pixel_row     : IN STD_LOGIC_VECTOR( 9 DOWNTO 0 );
	    o_red           : OUT STD_LOGIC_VECTOR( 7 DOWNTO 0 );
	    o_green         : OUT STD_LOGIC_VECTOR( 7 DOWNTO 0 );
	    o_blue          : OUT STD_LOGIC_VECTOR( 7 DOWNTO 0 ));
END color_rom_vhd; 

ARCHITECTURE behavioral OF color_rom_vhd  IS 

CONSTANT BATASBARIS   : INTEGER := 479;
CONSTANT BATASKOLOM   : INTEGER := 639;

SHARED VARIABLE LEVEL	: INTEGER := 1;
SHARED VARIABLE UTAMA	: BOOLEAN := FALSE;
SHARED VARIABLE MENANG	: BOOLEAN := FALSE;
SHARED VARIABLE KALAH	: BOOLEAN := FALSE;
SHARED VARIABLE	KALAH1	: BOOLEAN := FALSE;
SHARED VARIABLE RESTART	: BOOLEAN := FALSE;
SHARED VARIABLE RESET	: BOOLEAN := FALSE;

--AWAL LEVEL 1
SHARED VARIABLE B1_ATAS : INTEGER := 10; 
SHARED VARIABLE B1_KIRI : INTEGER := 10; 
SHARED VARIABLE B1_KANAN : INTEGER := 60; 
SHARED VARIABLE B1_BAWAH : INTEGER := 60; 

SHARED VARIABLE S_ATAS : INTEGER := 10; 
SHARED VARIABLE S_KIRI : INTEGER := 10; 
SHARED VARIABLE S_KANAN : INTEGER := 60; 
SHARED VARIABLE S_BAWAH : INTEGER := 60; 

SHARED VARIABLE GR1_ATAS : INTEGER := 0; 
SHARED VARIABLE GR1_KIRI : INTEGER := 0; 
SHARED VARIABLE GR1_KANAN : INTEGER := 10; 
SHARED VARIABLE GR1_BAWAH : INTEGER := 480;

SHARED VARIABLE GR2_ATAS : INTEGER := 0; 
SHARED VARIABLE GR2_KIRI : INTEGER := 0; 
SHARED VARIABLE GR2_KANAN : INTEGER := 639; 
SHARED VARIABLE GR2_BAWAH : INTEGER := 10; 

SHARED VARIABLE GR3_ATAS : INTEGER := 470; 
SHARED VARIABLE GR3_KIRI : INTEGER := 0; 
SHARED VARIABLE GR3_KANAN : INTEGER := 640; 
SHARED VARIABLE GR3_BAWAH : INTEGER := 480; 

SHARED VARIABLE GR4_ATAS : INTEGER := 0; 
SHARED VARIABLE GR4_KIRI : INTEGER := 620; 
SHARED VARIABLE GR4_KANAN : INTEGER := 630; 
SHARED VARIABLE GR4_BAWAH : INTEGER := 480;

SHARED VARIABLE GR5_ATAS : INTEGER := 140; 
SHARED VARIABLE GR5_KIRI : INTEGER := 0; 
SHARED VARIABLE GR5_KANAN : INTEGER := 140; 
SHARED VARIABLE GR5_BAWAH : INTEGER := 150;

SHARED VARIABLE GR6_ATAS : INTEGER := 210; 
SHARED VARIABLE GR6_KIRI : INTEGER := 0; 
SHARED VARIABLE GR6_KANAN : INTEGER := 140; 
SHARED VARIABLE GR6_BAWAH : INTEGER := 220;

SHARED VARIABLE GR8_ATAS : INTEGER := 340; 
SHARED VARIABLE GR8_KIRI : INTEGER := 70; 
SHARED VARIABLE GR8_KANAN : INTEGER := 140; 
SHARED VARIABLE GR8_BAWAH : INTEGER := 350;

SHARED VARIABLE GR9_ATAS : INTEGER := 410; 
SHARED VARIABLE GR9_KIRI : INTEGER := 130; 
SHARED VARIABLE GR9_KANAN : INTEGER := 330; 
SHARED VARIABLE GR9_BAWAH : INTEGER := 420;

SHARED VARIABLE GR10_ATAS : INTEGER := 280; 
SHARED VARIABLE GR10_KIRI : INTEGER := 190; 
SHARED VARIABLE GR10_KANAN : INTEGER := 420; 
SHARED VARIABLE GR10_BAWAH : INTEGER := 290;

SHARED VARIABLE GR11_ATAS : INTEGER := 90; 
SHARED VARIABLE GR11_KIRI : INTEGER := 300; 
SHARED VARIABLE GR11_KANAN : INTEGER := 380; 
SHARED VARIABLE GR11_BAWAH : INTEGER := 100;

SHARED VARIABLE GR12_ATAS : INTEGER := 90; 
SHARED VARIABLE GR12_KIRI : INTEGER := 470; 
SHARED VARIABLE GR12_KANAN : INTEGER := 570; 
SHARED VARIABLE GR12_BAWAH : INTEGER := 100;

SHARED VARIABLE GR13_ATAS : INTEGER := 310; 
SHARED VARIABLE GR13_KIRI : INTEGER := 470; 
SHARED VARIABLE GR13_KANAN : INTEGER := 570; 
SHARED VARIABLE GR13_BAWAH : INTEGER := 100;

SHARED VARIABLE GR14_ATAS : INTEGER := 400; 
SHARED VARIABLE GR14_KIRI : INTEGER := 560; 
SHARED VARIABLE GR14_KANAN : INTEGER := 630; 
SHARED VARIABLE GR14_BAWAH : INTEGER := 410;

SHARED VARIABLE GC1_ATAS  : INTEGER := 0; 
SHARED VARIABLE GC1_KIRI  : INTEGER := 80; 
SHARED VARIABLE GC1_KANAN : INTEGER := 90; 
SHARED VARIABLE GC1_BAWAH : INTEGER := 80;

SHARED VARIABLE GC2_ATAS  : INTEGER := 0; 
SHARED VARIABLE GC2_KIRI  : INTEGER := 220; 
SHARED VARIABLE GC2_KANAN : INTEGER := 230; 
SHARED VARIABLE GC2_BAWAH : INTEGER := 160;

SHARED VARIABLE GC3_ATAS  : INTEGER := 90; 
SHARED VARIABLE GC3_KIRI  : INTEGER := 360; 
SHARED VARIABLE GC3_KANAN : INTEGER := 370; 
SHARED VARIABLE GC3_BAWAH : INTEGER := 190;

SHARED VARIABLE GC4_ATAS  : INTEGER := 230; 
SHARED VARIABLE GC4_KIRI  : INTEGER := 270; 
SHARED VARIABLE GC4_KANAN : INTEGER := 280; 
SHARED VARIABLE GC4_BAWAH : INTEGER := 290;

SHARED VARIABLE GC5_ATAS  : INTEGER := 280; 
SHARED VARIABLE GC5_KIRI  : INTEGER := 60; 
SHARED VARIABLE GC5_KANAN : INTEGER := 70; 
SHARED VARIABLE GC5_BAWAH : INTEGER := 480;

SHARED VARIABLE GC7_ATAS  : INTEGER := 370; 
SHARED VARIABLE GC7_KIRI  : INTEGER := 400; 
SHARED VARIABLE GC7_KANAN : INTEGER := 410; 
SHARED VARIABLE GC7_BAWAH : INTEGER := 480;

SHARED VARIABLE GC8_ATAS  : INTEGER := 240; 
SHARED VARIABLE GC8_KIRI  : INTEGER := 460; 
SHARED VARIABLE GC8_KANAN : INTEGER := 470; 
SHARED VARIABLE GC8_BAWAH : INTEGER := 360;

SHARED VARIABLE F_ATAS : INTEGER := 410; 
SHARED VARIABLE F_KIRI : INTEGER := 570; 
SHARED VARIABLE F_KANAN : INTEGER := 630; 
SHARED VARIABLE F_BAWAH : INTEGER := 470;


--AWAL LEVEL 2
SHARED VARIABLE B_ATAS : INTEGER := 10; 
SHARED VARIABLE B_KIRI : INTEGER := 20; 
SHARED VARIABLE B_KANAN : INTEGER := 50; 
SHARED VARIABLE B_BAWAH : INTEGER := 40;

--PEMICU BATAS
SHARED VARIABLE P_ATAS : INTEGER := 10; 
SHARED VARIABLE P_KIRI : INTEGER := 20; 
SHARED VARIABLE P_KANAN : INTEGER := 50; 
SHARED VARIABLE P_BAWAH : INTEGER := 40; 

--BINGKAI ATAS
SHARED VARIABLE G1_ATAS : INTEGER := 0; 
SHARED VARIABLE G1_KIRI : INTEGER := 0; 
SHARED VARIABLE G1_KANAN : INTEGER := 640; 
SHARED VARIABLE G1_BAWAH : INTEGER := 10;

--BINGKAI KIRI
SHARED VARIABLE G2_ATAS : INTEGER := 0; 
SHARED VARIABLE G2_KIRI : INTEGER := 0; 
SHARED VARIABLE G2_KANAN : INTEGER := 10; 
SHARED VARIABLE G2_BAWAH : INTEGER := 480;

--BINGKAI BAWAH
SHARED VARIABLE G3_ATAS : INTEGER := 470; 
SHARED VARIABLE G3_KIRI : INTEGER := 0; 
SHARED VARIABLE G3_KANAN : INTEGER := 640; 
SHARED VARIABLE G3_BAWAH : INTEGER := 480;

--BINGKAI KANAN
SHARED VARIABLE G4_ATAS : INTEGER := 0; 
SHARED VARIABLE G4_KIRI : INTEGER := 620; 
SHARED VARIABLE G4_KANAN : INTEGER := 630; 
SHARED VARIABLE G4_BAWAH : INTEGER := 480;

--GARIS VERTIKAL ANTARA I DAN M
SHARED VARIABLE G5_ATAS : INTEGER := 0; 
SHARED VARIABLE G5_KIRI : INTEGER := 50; 
SHARED VARIABLE G5_KANAN : INTEGER := 60; 
SHARED VARIABLE G5_BAWAH : INTEGER := 170;

--GARIS HORIZONTAL I DAN M POJOK KIRI BAWAH
SHARED VARIABLE G6_ATAS : INTEGER := 160; 
SHARED VARIABLE G6_KIRI : INTEGER := 0; 
SHARED VARIABLE G6_KANAN : INTEGER := 110; 
SHARED VARIABLE G6_BAWAH : INTEGER := 170;

--GARIS VERTIKAL M_1
SHARED VARIABLE G7_ATAS : INTEGER := 50; 
SHARED VARIABLE G7_KIRI : INTEGER := 100; 
SHARED VARIABLE G7_KANAN : INTEGER := 110; 
SHARED VARIABLE G7_BAWAH : INTEGER := 170;

--GARIS VERTIKAL M_2 AMPE BAWAH
SHARED VARIABLE G8_ATAS : INTEGER := 50; 
SHARED VARIABLE G8_KIRI : INTEGER := 150; 
SHARED VARIABLE G8_KANAN : INTEGER := 160; 
SHARED VARIABLE G8_BAWAH : INTEGER := 480;

--GARIS VERTIKAL M_3
SHARED VARIABLE G9_ATAS : INTEGER := 50; 
SHARED VARIABLE G9_KIRI : INTEGER := 200; 
SHARED VARIABLE G9_KANAN : INTEGER := 210; 
SHARED VARIABLE G9_BAWAH : INTEGER := 170;

--GARIS VERTIKAL M_4
SHARED VARIABLE G10_ATAS : INTEGER := 50; 
SHARED VARIABLE G10_KIRI : INTEGER := 250; 
SHARED VARIABLE G10_KANAN : INTEGER := 260; 
SHARED VARIABLE G10_BAWAH : INTEGER := 170;

--GARIS HORIZONTAL M ATAS KIRI
SHARED VARIABLE G11_ATAS : INTEGER := 50; 
SHARED VARIABLE G11_KIRI : INTEGER := 100; 
SHARED VARIABLE G11_KANAN : INTEGER := 160; 
SHARED VARIABLE G11_BAWAH : INTEGER := 60;

--GARIS HORIZONTAL M ATAS KANAN
SHARED VARIABLE G12_ATAS : INTEGER := 50; 
SHARED VARIABLE G12_KIRI : INTEGER := 200; 
SHARED VARIABLE G12_KANAN : INTEGER := 260; 
SHARED VARIABLE G12_BAWAH : INTEGER := 60;

--GARIS HORIZONTAL M BAWAH
SHARED VARIABLE G13_ATAS : INTEGER := 160; 
SHARED VARIABLE G13_KIRI : INTEGER := 150; 
SHARED VARIABLE G13_KANAN : INTEGER := 210; 
SHARED VARIABLE G13_BAWAH : INTEGER := 170;

--GARIS HORIZONTAL M POJOK BAWAH KANAN AMPE A
SHARED VARIABLE G14_ATAS : INTEGER := 160; 
SHARED VARIABLE G14_KIRI : INTEGER := 250; 
SHARED VARIABLE G14_KANAN : INTEGER := 350; 
SHARED VARIABLE G14_BAWAH : INTEGER := 170;

--GARIS VERTIKAL ANTARA M DAN A
SHARED VARIABLE G15_ATAS : INTEGER := 0; 
SHARED VARIABLE G15_KIRI : INTEGER := 300; 
SHARED VARIABLE G15_KANAN : INTEGER := 310; 
SHARED VARIABLE G15_BAWAH : INTEGER := 170;

--KOTAK DI TENGAH A
SHARED VARIABLE G16_ATAS : INTEGER := 50; 
SHARED VARIABLE G16_KIRI : INTEGER := 350; 
SHARED VARIABLE G16_KANAN : INTEGER := 410; 
SHARED VARIABLE G16_BAWAH : INTEGER := 80;

--GARIS HORIZONTAL A TENGAH
SHARED VARIABLE G17_ATAS : INTEGER := 120; 
SHARED VARIABLE G17_KIRI : INTEGER := 350; 
SHARED VARIABLE G17_KANAN : INTEGER := 410; 
SHARED VARIABLE G17_BAWAH : INTEGER := 130;

--GARIS HORIZONTAL A POJOK KANAN BAWAH
SHARED VARIABLE G18_ATAS : INTEGER := 160; 
SHARED VARIABLE G18_KIRI : INTEGER := 400; 
SHARED VARIABLE G18_KANAN : INTEGER := 480; 
SHARED VARIABLE G18_BAWAH : INTEGER := 170;

--KOTAK DI KANAN A
SHARED VARIABLE G19_ATAS : INTEGER := 0; 
SHARED VARIABLE G19_KIRI : INTEGER := 450; 
SHARED VARIABLE G19_KANAN : INTEGER := 480; 
SHARED VARIABLE G19_BAWAH : INTEGER := 170;

--GARIS VERTIKAL A_1 AMPE UJUNG BAWAH
SHARED VARIABLE G20_ATAS : INTEGER := 120; 
SHARED VARIABLE G20_KIRI : INTEGER := 350; 
SHARED VARIABLE G20_KANAN : INTEGER := 360; 
SHARED VARIABLE G20_BAWAH : INTEGER := 480;

--GARIS VERTIKAL A_2 AMPE LEKUKAN BAWAH
SHARED VARIABLE G21_ATAS : INTEGER := 120; 
SHARED VARIABLE G21_KIRI : INTEGER := 400; 
SHARED VARIABLE G21_KANAN : INTEGER := 410; 
SHARED VARIABLE G21_BAWAH : INTEGER := 430;

--KOTAK DI BAWAH I
SHARED VARIABLE G22_ATAS : INTEGER := 160; 
SHARED VARIABLE G22_KIRI : INTEGER := 50; 
SHARED VARIABLE G22_KANAN : INTEGER := 110; 
SHARED VARIABLE G22_BAWAH : INTEGER := 280;

--GARIS HORIZONTAL_1 DI BAWAH I
SHARED VARIABLE G23_ATAS : INTEGER := 320; 
SHARED VARIABLE G23_KIRI : INTEGER := 0; 
SHARED VARIABLE G23_KANAN : INTEGER := 110; 
SHARED VARIABLE G23_BAWAH : INTEGER := 330;

--GARIS HORIZONTAL_2 DI BAWAH I
SHARED VARIABLE G24_ATAS : INTEGER := 370; 
SHARED VARIABLE G24_KIRI : INTEGER := 0; 
SHARED VARIABLE G24_KANAN : INTEGER := 160; 
SHARED VARIABLE G24_BAWAH : INTEGER := 380;

--GARIS HORIZONTAL_3 DI BAWAH I
SHARED VARIABLE G25_ATAS : INTEGER := 420; 
SHARED VARIABLE G25_KIRI : INTEGER := 0; 
SHARED VARIABLE G25_KANAN : INTEGER := 110; 
SHARED VARIABLE G25_BAWAH : INTEGER := 430;

--GARIS HORIZONTAL_1 DI BAWAH M
SHARED VARIABLE G26_ATAS : INTEGER := 220; 
SHARED VARIABLE G26_KIRI : INTEGER := 200; 
SHARED VARIABLE G26_KANAN : INTEGER := 360; 
SHARED VARIABLE G26_BAWAH : INTEGER := 230;

--KOTAK DIBAWAH M
SHARED VARIABLE G27_ATAS : INTEGER := 270; 
SHARED VARIABLE G27_KIRI : INTEGER := 200; 
SHARED VARIABLE G27_KANAN : INTEGER := 310; 
SHARED VARIABLE G27_BAWAH : INTEGER := 320;

--GARIS VERTIKAL_1 DI BAWAH M
SHARED VARIABLE G28_ATAS : INTEGER := 270; 
SHARED VARIABLE G28_KIRI : INTEGER := 200; 
SHARED VARIABLE G28_KANAN : INTEGER := 210; 
SHARED VARIABLE G28_BAWAH : INTEGER := 370;

--GARIS VERTIKAL_2 DI BAWAH M
SHARED VARIABLE G29_ATAS : INTEGER := 270; 
SHARED VARIABLE G29_KIRI : INTEGER := 300; 
SHARED VARIABLE G29_KANAN : INTEGER := 310; 
SHARED VARIABLE G29_BAWAH : INTEGER := 340;

--GARIS HORIZONTAL_2 DI BAWAH M
SHARED VARIABLE G30_ATAS : INTEGER := 360; 
SHARED VARIABLE G30_KIRI : INTEGER := 200; 
SHARED VARIABLE G30_KANAN : INTEGER := 310; 
SHARED VARIABLE G30_BAWAH : INTEGER := 370;

--GARIS HORIZONTAL_3 DI BAWAH M
SHARED VARIABLE G31_ATAS : INTEGER := 420; 
SHARED VARIABLE G31_KIRI : INTEGER := 200; 
SHARED VARIABLE G31_KANAN : INTEGER := 360; 
SHARED VARIABLE G31_BAWAH : INTEGER := 430;

--GARIS HORIZONTAL DI BAWAH A
SHARED VARIABLE G32_ATAS : INTEGER := 420; 
SHARED VARIABLE G32_KIRI : INTEGER := 400; 
SHARED VARIABLE G32_KANAN : INTEGER := 450; 
SHARED VARIABLE G32_BAWAH : INTEGER := 430;

--KOTAK DI BAWAH A
SHARED VARIABLE G33_ATAS : INTEGER := 210; 
SHARED VARIABLE G33_KIRI : INTEGER := 450; 
SHARED VARIABLE G33_KANAN : INTEGER := 500; 
SHARED VARIABLE G33_BAWAH : INTEGER := 370;

--GARIS VERTIKAL DI BAWAH A
SHARED VARIABLE G34_ATAS : INTEGER := 210; 
SHARED VARIABLE G34_KIRI : INTEGER := 490; 
SHARED VARIABLE G34_KANAN : INTEGER := 500; 
SHARED VARIABLE G34_BAWAH : INTEGER := 480;

--GARIS VERTIKAL_1 DI KANAN A
SHARED VARIABLE G35_ATAS : INTEGER := 0; 
SHARED VARIABLE G35_KIRI : INTEGER := 520; 
SHARED VARIABLE G35_KANAN : INTEGER := 530; 
SHARED VARIABLE G35_BAWAH : INTEGER := 140;

--GARIS VERTIKAL_2 DI KANAN A
SHARED VARIABLE G36_ATAS : INTEGER := 0; 
SHARED VARIABLE G36_KIRI : INTEGER := 570; 
SHARED VARIABLE G36_KANAN : INTEGER := 580; 
SHARED VARIABLE G36_BAWAH : INTEGER := 190;

--GARIS HORIZONTAL DI KANAN A
SHARED VARIABLE G37_ATAS : INTEGER := 130; 
SHARED VARIABLE G37_KIRI : INTEGER := 520; 
SHARED VARIABLE G37_KANAN : INTEGER := 580; 
SHARED VARIABLE G37_BAWAH : INTEGER := 140;

--GARIS VERTIKAL_1 DI BAWAH U
SHARED VARIABLE G40_ATAS : INTEGER := 180; 
SHARED VARIABLE G40_KIRI : INTEGER := 540; 
SHARED VARIABLE G40_KANAN : INTEGER := 550; 
SHARED VARIABLE G40_BAWAH : INTEGER := 420;

--GARIS VERTIKAL_2 DI BAWAH U
SHARED VARIABLE G41_ATAS : INTEGER := 220; 
SHARED VARIABLE G41_KIRI : INTEGER := 580; 
SHARED VARIABLE G41_KANAN : INTEGER := 590; 
SHARED VARIABLE G41_BAWAH : INTEGER := 260;

--GARIS HORIZONTAL_1 DI BAWAH U
SHARED VARIABLE G42_ATAS : INTEGER := 180; 
SHARED VARIABLE G42_KIRI : INTEGER := 540; 
SHARED VARIABLE G42_KANAN : INTEGER := 630; 
SHARED VARIABLE G42_BAWAH : INTEGER := 190;

--GARIS HORIZONTAL_3 DI BAWAH U
SHARED VARIABLE G44_ATAS : INTEGER := 310; 
SHARED VARIABLE G44_KIRI : INTEGER := 540; 
SHARED VARIABLE G44_KANAN : INTEGER := 590; 
SHARED VARIABLE G44_BAWAH : INTEGER := 320;

--GARIS HORIZONTAL_4 DI BAWAH U
SHARED VARIABLE G45_ATAS : INTEGER := 360; 
SHARED VARIABLE G45_KIRI : INTEGER := 580; 
SHARED VARIABLE G45_KANAN : INTEGER := 630; 
SHARED VARIABLE G45_BAWAH : INTEGER := 370;

--GARIS HORIZONTAL_5 DI BAWAH U
SHARED VARIABLE G46_ATAS : INTEGER := 410; 
SHARED VARIABLE G46_KIRI : INTEGER := 540; 
SHARED VARIABLE G46_KANAN : INTEGER := 590; 
SHARED VARIABLE G46_BAWAH : INTEGER := 420;

--TELEPORT 1
SHARED VARIABLE G47_ATAS : INTEGER := 120; 
SHARED VARIABLE G47_KIRI : INTEGER := 10; 
SHARED VARIABLE G47_KANAN : INTEGER := 50; 
SHARED VARIABLE G47_BAWAH : INTEGER := 160;

--TELEPORT 2
SHARED VARIABLE G48_ATAS : INTEGER := 120; 
SHARED VARIABLE G48_KIRI : INTEGER := 60; 
SHARED VARIABLE G48_KANAN : INTEGER := 100; 
SHARED VARIABLE G48_BAWAH : INTEGER := 160;

--TELEPORT 3
SHARED VARIABLE G49_ATAS : INTEGER := 60; 
SHARED VARIABLE G49_KIRI : INTEGER := 110; 
SHARED VARIABLE G49_KANAN : INTEGER := 150; 
SHARED VARIABLE G49_BAWAH : INTEGER := 100;

--TELEPORT 4
SHARED VARIABLE G50_ATAS : INTEGER := 120; 
SHARED VARIABLE G50_KIRI : INTEGER := 260; 
SHARED VARIABLE G50_KANAN : INTEGER := 300; 
SHARED VARIABLE G50_BAWAH : INTEGER := 160;

--TELEPORT 5
SHARED VARIABLE G51_ATAS : INTEGER := 120; 
SHARED VARIABLE G51_KIRI : INTEGER := 310; 
SHARED VARIABLE G51_KANAN : INTEGER := 350; 
SHARED VARIABLE G51_BAWAH : INTEGER := 160;

--TELEPORT 6
SHARED VARIABLE G52_ATAS : INTEGER := 120; 
SHARED VARIABLE G52_KIRI : INTEGER := 410; 
SHARED VARIABLE G52_KANAN : INTEGER := 450; 
SHARED VARIABLE G52_BAWAH : INTEGER := 160;

--TELEPORT 7
SHARED VARIABLE G53_ATAS : INTEGER := 330; 
SHARED VARIABLE G53_KIRI : INTEGER := 10; 
SHARED VARIABLE G53_KANAN : INTEGER := 50; 
SHARED VARIABLE G53_BAWAH : INTEGER := 370;

--TELEPORT 8
SHARED VARIABLE G54_ATAS : INTEGER := 430; 
SHARED VARIABLE G54_KIRI : INTEGER := 10; 
SHARED VARIABLE G54_KANAN : INTEGER := 50; 
SHARED VARIABLE G54_BAWAH : INTEGER := 470;

--TELEPORT 9
SHARED VARIABLE G55_ATAS : INTEGER := 320; 
SHARED VARIABLE G55_KIRI : INTEGER := 210; 
SHARED VARIABLE G55_KANAN : INTEGER := 250; 
SHARED VARIABLE G55_BAWAH : INTEGER := 360;

--TELEPORT 10
SHARED VARIABLE G56_ATAS : INTEGER := 430; 
SHARED VARIABLE G56_KIRI : INTEGER := 310; 
SHARED VARIABLE G56_KANAN : INTEGER := 350; 
SHARED VARIABLE G56_BAWAH : INTEGER := 470;

--TELEPORT 11
SHARED VARIABLE G57_ATAS : INTEGER := 10; 
SHARED VARIABLE G57_KIRI : INTEGER := 530; 
SHARED VARIABLE G57_KANAN : INTEGER := 570; 
SHARED VARIABLE G57_BAWAH : INTEGER := 50;

--TELEPORT 12
SHARED VARIABLE G58_ATAS : INTEGER := 220; 
SHARED VARIABLE G58_KIRI : INTEGER := 590; 
SHARED VARIABLE G58_KANAN : INTEGER := 620; 
SHARED VARIABLE G58_BAWAH : INTEGER := 260;

--TELEPORT 13
SHARED VARIABLE G59_ATAS : INTEGER := 190; 
SHARED VARIABLE G59_KIRI : INTEGER := 590; 
SHARED VARIABLE G59_KANAN : INTEGER := 620; 
SHARED VARIABLE G59_BAWAH : INTEGER := 230;

--TELEPORT 14
SHARED VARIABLE G60_ATAS : INTEGER := 60; 
SHARED VARIABLE G60_KIRI : INTEGER := 210; 
SHARED VARIABLE G60_KANAN : INTEGER := 250; 
SHARED VARIABLE G60_BAWAH : INTEGER := 100;

--FINISH
SHARED VARIABLE G61_ATAS : INTEGER := 10; 
SHARED VARIABLE G61_KIRI : INTEGER := 580; 
SHARED VARIABLE G61_KANAN : INTEGER := 620; 
SHARED VARIABLE G61_BAWAH : INTEGER := 50;

--WAKTU LEVEL 1
SHARED VARIABLE G62_ATAS : INTEGER := 10; 
SHARED VARIABLE G62_KIRI : INTEGER := 630; 
SHARED VARIABLE G62_KANAN : INTEGER := 640; 
SHARED VARIABLE G62_BAWAH : INTEGER := 470;

SHARED VARIABLE G62A_ATAS : INTEGER := 10; 
SHARED VARIABLE G62A_KIRI : INTEGER := 630; 
SHARED VARIABLE G62A_KANAN : INTEGER := 640; 
SHARED VARIABLE G62A_BAWAH : INTEGER := 470;

SHARED VARIABLE G62B_ATAS : INTEGER := 10; 
SHARED VARIABLE G62B_KIRI : INTEGER := 630; 
SHARED VARIABLE G62B_KANAN : INTEGER := 640; 
SHARED VARIABLE G62B_BAWAH : INTEGER := 470;

--WAKTU LEVEL 2
SHARED VARIABLE G63_ATAS : INTEGER := 10; 
SHARED VARIABLE G63_KIRI : INTEGER := 630; 
SHARED VARIABLE G63_KANAN : INTEGER := 640; 
SHARED VARIABLE G63_BAWAH : INTEGER := 470;

SHARED VARIABLE G63A_ATAS : INTEGER := 10; 
SHARED VARIABLE G63A_KIRI : INTEGER := 630; 
SHARED VARIABLE G63A_KANAN : INTEGER := 640; 
SHARED VARIABLE G63A_BAWAH : INTEGER := 470;

SHARED VARIABLE G63B_ATAS : INTEGER := 10; 
SHARED VARIABLE G63B_KIRI : INTEGER := 630; 
SHARED VARIABLE G63B_KANAN : INTEGER := 640; 
SHARED VARIABLE G63B_BAWAH : INTEGER := 470;


--LAYAR AWAL

--HURUF I
SHARED VARIABLE G64_ATAS : INTEGER := 120; 
SHARED VARIABLE G64_KIRI : INTEGER := 200; 
SHARED VARIABLE G64_KANAN : INTEGER := 210; 
SHARED VARIABLE G64_BAWAH : INTEGER := 250;

--GARIS M KIRI
SHARED VARIABLE G65_ATAS : INTEGER := 120; 
SHARED VARIABLE G65_KIRI : INTEGER := 230; 
SHARED VARIABLE G65_KANAN : INTEGER := 240; 
SHARED VARIABLE G65_BAWAH : INTEGER := 250;

--GARIS M TENGAH
SHARED VARIABLE G66_ATAS : INTEGER := 120; 
SHARED VARIABLE G66_KIRI : INTEGER := 280; 
SHARED VARIABLE G66_KANAN : INTEGER := 290; 
SHARED VARIABLE G66_BAWAH : INTEGER := 250;

--GARIS M KANAN
SHARED VARIABLE G67_ATAS : INTEGER := 120; 
SHARED VARIABLE G67_KIRI : INTEGER := 330; 
SHARED VARIABLE G67_KANAN : INTEGER := 340; 
SHARED VARIABLE G67_BAWAH : INTEGER := 250;

--GARIS M ATAS
SHARED VARIABLE G68_ATAS : INTEGER := 120; 
SHARED VARIABLE G68_KIRI : INTEGER := 230; 
SHARED VARIABLE G68_KANAN : INTEGER := 340; 
SHARED VARIABLE G68_BAWAH : INTEGER := 130;

--GARIS KIRI A
SHARED VARIABLE G69_ATAS : INTEGER := 120; 
SHARED VARIABLE G69_KIRI : INTEGER := 360; 
SHARED VARIABLE G69_KANAN : INTEGER := 370; 
SHARED VARIABLE G69_BAWAH : INTEGER := 250;

--GARIS KANAN A
SHARED VARIABLE G70_ATAS : INTEGER := 120; 
SHARED VARIABLE G70_KIRI : INTEGER := 420; 
SHARED VARIABLE G70_KANAN : INTEGER := 430; 
SHARED VARIABLE G70_BAWAH : INTEGER := 250;

--GARIS ATAS A
SHARED VARIABLE G71_ATAS : INTEGER := 120; 
SHARED VARIABLE G71_KIRI : INTEGER := 360; 
SHARED VARIABLE G71_KANAN : INTEGER := 430; 
SHARED VARIABLE G71_BAWAH : INTEGER := 130;

--GARIS TENGAH A
SHARED VARIABLE G72_ATAS : INTEGER := 180; 
SHARED VARIABLE G72_KIRI : INTEGER := 360; 
SHARED VARIABLE G72_KANAN : INTEGER := 430; 
SHARED VARIABLE G72_BAWAH : INTEGER := 190;

--GARIS L_1
SHARED VARIABLE G73_ATAS : INTEGER := 280; 
SHARED VARIABLE G73_KIRI : INTEGER := 170; 
SHARED VARIABLE G73_KANAN : INTEGER := 180; 
SHARED VARIABLE G73_BAWAH : INTEGER := 330;

--GARIS L_2
SHARED VARIABLE G74_ATAS : INTEGER := 320; 
SHARED VARIABLE G74_KIRI : INTEGER := 170; 
SHARED VARIABLE G74_KANAN : INTEGER := 210; 
SHARED VARIABLE G74_BAWAH : INTEGER := 330;

--GARIS E_1
SHARED VARIABLE G75_ATAS : INTEGER := 280; 
SHARED VARIABLE G75_KIRI : INTEGER := 220; 
SHARED VARIABLE G75_KANAN : INTEGER := 230; 
SHARED VARIABLE G75_BAWAH : INTEGER := 330;

--GARIS E_2
SHARED VARIABLE G76_ATAS : INTEGER := 280; 
SHARED VARIABLE G76_KIRI : INTEGER := 220; 
SHARED VARIABLE G76_KANAN : INTEGER := 260; 
SHARED VARIABLE G76_BAWAH : INTEGER := 290;

--GARIS E_3
SHARED VARIABLE G77_ATAS : INTEGER := 300; 
SHARED VARIABLE G77_KIRI : INTEGER := 220; 
SHARED VARIABLE G77_KANAN : INTEGER := 260; 
SHARED VARIABLE G77_BAWAH : INTEGER := 310;

--GARIS E_4
SHARED VARIABLE G78_ATAS : INTEGER := 320; 
SHARED VARIABLE G78_KIRI : INTEGER := 220; 
SHARED VARIABLE G78_KANAN : INTEGER := 260; 
SHARED VARIABLE G78_BAWAH : INTEGER := 330;

--GARIS G_1
SHARED VARIABLE G79_ATAS : INTEGER := 280; 
SHARED VARIABLE G79_KIRI : INTEGER := 270; 
SHARED VARIABLE G79_KANAN : INTEGER := 280; 
SHARED VARIABLE G79_BAWAH : INTEGER := 330;

--GARIS G_2
SHARED VARIABLE G80_ATAS : INTEGER := 300; 
SHARED VARIABLE G80_KIRI : INTEGER := 300; 
SHARED VARIABLE G80_KANAN : INTEGER := 310; 
SHARED VARIABLE G80_BAWAH : INTEGER := 330;

--GARIS G_3
SHARED VARIABLE G81_ATAS : INTEGER := 280; 
SHARED VARIABLE G81_KIRI : INTEGER := 270; 
SHARED VARIABLE G81_KANAN : INTEGER := 310; 
SHARED VARIABLE G81_BAWAH : INTEGER := 290;

--GARIS G_4
SHARED VARIABLE G82_ATAS : INTEGER := 300; 
SHARED VARIABLE G82_KIRI : INTEGER := 290; 
SHARED VARIABLE G82_KANAN : INTEGER := 310; 
SHARED VARIABLE G82_BAWAH : INTEGER := 310;

--GARIS G_5
SHARED VARIABLE G83_ATAS : INTEGER := 320; 
SHARED VARIABLE G83_KIRI : INTEGER := 270; 
SHARED VARIABLE G83_KANAN : INTEGER := 310; 
SHARED VARIABLE G83_BAWAH : INTEGER := 330;

--GARIS E_5
SHARED VARIABLE G84_ATAS : INTEGER := 280; 
SHARED VARIABLE G84_KIRI : INTEGER := 320; 
SHARED VARIABLE G84_KANAN : INTEGER := 330; 
SHARED VARIABLE G84_BAWAH : INTEGER := 330;

--GARIS E_6
SHARED VARIABLE G85_ATAS : INTEGER := 280; 
SHARED VARIABLE G85_KIRI : INTEGER := 320; 
SHARED VARIABLE G85_KANAN : INTEGER := 360; 
SHARED VARIABLE G85_BAWAH : INTEGER := 290;

--GARIS E_7
SHARED VARIABLE G86_ATAS : INTEGER := 300; 
SHARED VARIABLE G86_KIRI : INTEGER := 320; 
SHARED VARIABLE G86_KANAN : INTEGER := 360; 
SHARED VARIABLE G86_BAWAH : INTEGER := 310;

--GARIS E_8
SHARED VARIABLE G87_ATAS : INTEGER := 320; 
SHARED VARIABLE G87_KIRI : INTEGER := 320; 
SHARED VARIABLE G87_KANAN : INTEGER := 360; 
SHARED VARIABLE G87_BAWAH : INTEGER := 330;

--GARIS N_1
SHARED VARIABLE G88_ATAS : INTEGER := 280; 
SHARED VARIABLE G88_KIRI : INTEGER := 370; 
SHARED VARIABLE G88_KANAN : INTEGER := 380; 
SHARED VARIABLE G88_BAWAH : INTEGER := 330;

--GARIS N_2
SHARED VARIABLE G89_ATAS : INTEGER := 280; 
SHARED VARIABLE G89_KIRI : INTEGER := 400; 
SHARED VARIABLE G89_KANAN : INTEGER := 410; 
SHARED VARIABLE G89_BAWAH : INTEGER := 330;

--GARIS N_3
SHARED VARIABLE G90_ATAS : INTEGER := 290; 
SHARED VARIABLE G90_KIRI : INTEGER := 370; 
SHARED VARIABLE G90_KANAN : INTEGER := 390; 
SHARED VARIABLE G90_BAWAH : INTEGER := 300;

--GARIS N_4
SHARED VARIABLE G91_ATAS : INTEGER := 310; 
SHARED VARIABLE G91_KIRI : INTEGER := 390; 
SHARED VARIABLE G91_KANAN : INTEGER := 410; 
SHARED VARIABLE G91_BAWAH : INTEGER := 320;

--GARIS D_1
SHARED VARIABLE G92_ATAS : INTEGER := 280; 
SHARED VARIABLE G92_KIRI : INTEGER := 420; 
SHARED VARIABLE G92_KANAN : INTEGER := 430; 
SHARED VARIABLE G92_BAWAH : INTEGER := 330;

--GARIS D_2
SHARED VARIABLE G93_ATAS : INTEGER := 290; 
SHARED VARIABLE G93_KIRI : INTEGER := 450; 
SHARED VARIABLE G93_KANAN : INTEGER := 460; 
SHARED VARIABLE G93_BAWAH : INTEGER := 320;

--GARIS D_3
SHARED VARIABLE G94_ATAS : INTEGER := 280; 
SHARED VARIABLE G94_KIRI : INTEGER := 420; 
SHARED VARIABLE G94_KANAN : INTEGER := 450; 
SHARED VARIABLE G94_BAWAH : INTEGER := 290;

--GARIS D_4
SHARED VARIABLE G95_ATAS : INTEGER := 320; 
SHARED VARIABLE G95_KIRI : INTEGER := 420; 
SHARED VARIABLE G95_KANAN : INTEGER := 450; 
SHARED VARIABLE G95_BAWAH : INTEGER := 330;

--GARIS Y_1
SHARED VARIABLE G96_ATAS : INTEGER := 390; 
SHARED VARIABLE G96_KIRI : INTEGER := 270; 
SHARED VARIABLE G96_KANAN : INTEGER := 280; 
SHARED VARIABLE G96_BAWAH : INTEGER := 410;

--GARIS Y_2
SHARED VARIABLE G97_ATAS : INTEGER := 390; 
SHARED VARIABLE G97_KIRI : INTEGER := 300; 
SHARED VARIABLE G97_KANAN : INTEGER := 310; 
SHARED VARIABLE G97_BAWAH : INTEGER := 410;

--GARIS Y_3
SHARED VARIABLE G98_ATAS : INTEGER := 410; 
SHARED VARIABLE G98_KIRI : INTEGER := 280; 
SHARED VARIABLE G98_KANAN : INTEGER := 300; 
SHARED VARIABLE G98_BAWAH : INTEGER := 420;

--GARIS Y_4
SHARED VARIABLE G99_ATAS : INTEGER := 410; 
SHARED VARIABLE G99_KIRI : INTEGER := 285; 
SHARED VARIABLE G99_KANAN : INTEGER := 295; 
SHARED VARIABLE G99_BAWAH : INTEGER := 440;

--GARIS 5_1
SHARED VARIABLE G100_ATAS : INTEGER := 390; 
SHARED VARIABLE G100_KIRI : INTEGER := 320; 
SHARED VARIABLE G100_KANAN : INTEGER := 360; 
SHARED VARIABLE G100_BAWAH : INTEGER := 400;

--GARIS 5_2
SHARED VARIABLE G101_ATAS : INTEGER := 410; 
SHARED VARIABLE G101_KIRI : INTEGER := 320; 
SHARED VARIABLE G101_KANAN : INTEGER := 360; 
SHARED VARIABLE G101_BAWAH : INTEGER := 420;

--GARIS 5_3
SHARED VARIABLE G102_ATAS : INTEGER := 430; 
SHARED VARIABLE G102_KIRI : INTEGER := 320; 
SHARED VARIABLE G102_KANAN : INTEGER := 360; 
SHARED VARIABLE G102_BAWAH : INTEGER := 440;

--GARIS 5_4
SHARED VARIABLE G103_ATAS : INTEGER := 390; 
SHARED VARIABLE G103_KIRI : INTEGER := 320; 
SHARED VARIABLE G103_KANAN : INTEGER := 330; 
SHARED VARIABLE G103_BAWAH : INTEGER := 420;

--GARIS 5_5
SHARED VARIABLE G104_ATAS : INTEGER := 410; 
SHARED VARIABLE G104_KIRI : INTEGER := 350; 
SHARED VARIABLE G104_KANAN : INTEGER := 360; 
SHARED VARIABLE G104_BAWAH : INTEGER := 440;


--KALAH

--GARIS L_1
SHARED VARIABLE G105_ATAS : INTEGER := 70; 
SHARED VARIABLE G105_KIRI : INTEGER := 110; 
SHARED VARIABLE G105_KANAN : INTEGER := 120; 
SHARED VARIABLE G105_BAWAH : INTEGER := 380;

--GARIS L_2
SHARED VARIABLE G106_ATAS : INTEGER := 370; 
SHARED VARIABLE G106_KIRI : INTEGER := 110; 
SHARED VARIABLE G106_KANAN : INTEGER := 190; 
SHARED VARIABLE G106_BAWAH : INTEGER := 380;

--GARIS O_1
SHARED VARIABLE G107_ATAS : INTEGER := 70; 
SHARED VARIABLE G107_KIRI : INTEGER := 220; 
SHARED VARIABLE G107_KANAN : INTEGER := 230; 
SHARED VARIABLE G107_BAWAH : INTEGER := 380;

--GARIS O_2
SHARED VARIABLE G108_ATAS : INTEGER := 70; 
SHARED VARIABLE G108_KIRI : INTEGER := 290; 
SHARED VARIABLE G108_KANAN : INTEGER := 300; 
SHARED VARIABLE G108_BAWAH : INTEGER := 380;

--GARIS O_3
SHARED VARIABLE G109_ATAS : INTEGER := 70; 
SHARED VARIABLE G109_KIRI : INTEGER := 220; 
SHARED VARIABLE G109_KANAN : INTEGER := 300; 
SHARED VARIABLE G109_BAWAH : INTEGER := 80;

--GARIS 0_4
SHARED VARIABLE G110_ATAS : INTEGER := 370; 
SHARED VARIABLE G110_KIRI : INTEGER := 220; 
SHARED VARIABLE G110_KANAN : INTEGER := 300; 
SHARED VARIABLE G110_BAWAH : INTEGER := 380;

--GARIS S_1
SHARED VARIABLE G111_ATAS : INTEGER := 70; 
SHARED VARIABLE G111_KIRI : INTEGER := 330; 
SHARED VARIABLE G111_KANAN : INTEGER := 340; 
SHARED VARIABLE G111_BAWAH : INTEGER := 220;

--GARIS S_2
SHARED VARIABLE G112_ATAS : INTEGER := 210; 
SHARED VARIABLE G112_KIRI : INTEGER := 400; 
SHARED VARIABLE G112_KANAN : INTEGER := 410; 
SHARED VARIABLE G112_BAWAH : INTEGER := 380;

--GARIS S_3
SHARED VARIABLE G113_ATAS : INTEGER := 70; 
SHARED VARIABLE G113_KIRI : INTEGER := 330; 
SHARED VARIABLE G113_KANAN : INTEGER := 410; 
SHARED VARIABLE G113_BAWAH : INTEGER := 80;

--GARIS S_4
SHARED VARIABLE G114_ATAS : INTEGER := 210; 
SHARED VARIABLE G114_KIRI : INTEGER := 330; 
SHARED VARIABLE G114_KANAN : INTEGER := 410; 
SHARED VARIABLE G114_BAWAH : INTEGER := 220;

--GARIS S_5
SHARED VARIABLE G115_ATAS : INTEGER := 370; 
SHARED VARIABLE G115_KIRI : INTEGER := 330; 
SHARED VARIABLE G115_KANAN : INTEGER := 410; 
SHARED VARIABLE G115_BAWAH : INTEGER := 380;

--GARIS E_1
SHARED VARIABLE G116_ATAS : INTEGER := 70; 
SHARED VARIABLE G116_KIRI : INTEGER := 440; 
SHARED VARIABLE G116_KANAN : INTEGER := 450; 
SHARED VARIABLE G116_BAWAH : INTEGER := 380;

--GARIS E_2
SHARED VARIABLE G117_ATAS : INTEGER := 70; 
SHARED VARIABLE G117_KIRI : INTEGER := 440; 
SHARED VARIABLE G117_KANAN : INTEGER := 520; 
SHARED VARIABLE G117_BAWAH : INTEGER := 80;

--GARIS E_3
SHARED VARIABLE G118_ATAS : INTEGER := 220; 
SHARED VARIABLE G118_KIRI : INTEGER := 440; 
SHARED VARIABLE G118_KANAN : INTEGER := 520; 
SHARED VARIABLE G118_BAWAH : INTEGER := 230;

--GARIS E_4
SHARED VARIABLE G119_ATAS : INTEGER := 370; 
SHARED VARIABLE G119_KIRI : INTEGER := 440; 
SHARED VARIABLE G119_KANAN : INTEGER := 520; 
SHARED VARIABLE G119_BAWAH : INTEGER := 380;


--MENANG

--GARIS W_1
SHARED VARIABLE G120_ATAS : INTEGER := 70; 
SHARED VARIABLE G120_KIRI : INTEGER := 150; 
SHARED VARIABLE G120_KANAN : INTEGER := 160; 
SHARED VARIABLE G120_BAWAH : INTEGER := 380;

--GARIS W_2
SHARED VARIABLE G121_ATAS : INTEGER := 70; 
SHARED VARIABLE G121_KIRI : INTEGER := 210; 
SHARED VARIABLE G121_KANAN : INTEGER := 220; 
SHARED VARIABLE G121_BAWAH : INTEGER := 380;

--GARIS W_3
SHARED VARIABLE G122_ATAS : INTEGER := 70; 
SHARED VARIABLE G122_KIRI : INTEGER := 270; 
SHARED VARIABLE G122_KANAN : INTEGER := 280; 
SHARED VARIABLE G122_BAWAH : INTEGER := 380;

--GARIS W_4
SHARED VARIABLE G123_ATAS : INTEGER := 370; 
SHARED VARIABLE G123_KIRI : INTEGER := 150; 
SHARED VARIABLE G123_KANAN : INTEGER := 280; 
SHARED VARIABLE G123_BAWAH : INTEGER := 380;

--GARIS I
SHARED VARIABLE G124_ATAS : INTEGER := 70; 
SHARED VARIABLE G124_KIRI : INTEGER := 310; 
SHARED VARIABLE G124_KANAN : INTEGER := 320; 
SHARED VARIABLE G124_BAWAH : INTEGER := 380;

--GARIS N_1
SHARED VARIABLE G125_ATAS : INTEGER := 70; 
SHARED VARIABLE G125_KIRI : INTEGER := 350; 
SHARED VARIABLE G125_KANAN : INTEGER := 360; 
SHARED VARIABLE G125_BAWAH : INTEGER := 380;

--GARIS N_2
SHARED VARIABLE G126_ATAS : INTEGER := 80; 
SHARED VARIABLE G126_KIRI : INTEGER := 400; 
SHARED VARIABLE G126_KANAN : INTEGER := 410; 
SHARED VARIABLE G126_BAWAH : INTEGER := 210;

--GARIS N_3
SHARED VARIABLE G127_ATAS : INTEGER := 210; 
SHARED VARIABLE G127_KIRI : INTEGER := 410; 
SHARED VARIABLE G127_KANAN : INTEGER := 420; 
SHARED VARIABLE G127_BAWAH : INTEGER := 240;

--GARIS N_4
SHARED VARIABLE G128_ATAS : INTEGER := 240; 
SHARED VARIABLE G128_KIRI : INTEGER := 420; 
SHARED VARIABLE G128_KANAN : INTEGER := 430; 
SHARED VARIABLE G128_BAWAH : INTEGER := 380;

--GARIS N_5
SHARED VARIABLE G129_ATAS : INTEGER := 70; 
SHARED VARIABLE G129_KIRI : INTEGER := 470; 
SHARED VARIABLE G129_KANAN : INTEGER := 480; 
SHARED VARIABLE G129_BAWAH : INTEGER := 380;

--GARIS N_6
SHARED VARIABLE G130_ATAS : INTEGER := 70; 
SHARED VARIABLE G130_KIRI : INTEGER := 350; 
SHARED VARIABLE G130_KANAN : INTEGER := 400; 
SHARED VARIABLE G130_BAWAH : INTEGER := 80;

--GARIS N_7
SHARED VARIABLE G131_ATAS : INTEGER := 370; 
SHARED VARIABLE G131_KIRI : INTEGER := 430; 
SHARED VARIABLE G131_KANAN : INTEGER := 480; 
SHARED VARIABLE G131_BAWAH : INTEGER := 380;

SIGNAL M_TF1, M_TF2                 :  STD_LOGIC; 
SIGNAL K_TF1, K_TF2                 :  STD_LOGIC; 
SIGNAL H_TF1, H_TF2                 :  STD_LOGIC; 

SHARED VARIABLE KECEPATAN 	: INTEGER 		:= 0;
SHARED VARIABLE KECEPATAN1	: INTEGER		:= 0;
SIGNAL clock40hz : STD_LOGIC;

COMPONENT CLOCKDIV is 
	port ( CLK : IN std_logic;
			DIVOUT : buffer std_logic);
end component;		

BEGIN 

PROCESS(i_pixel_row,i_pixel_column, i_M_US  , 
i_K_US  , i_H_US  , i_M_BT  , i_K_BT  , i_H_BT,
 M_TF1, M_TF2, K_TF1, K_TF2, H_TF1, H_TF2)

BEGIN

--LAYAR UTAMA
IF UTAMA = TRUE THEN
	IF ((i_pixel_column > G64_KIRI) AND (i_pixel_column < G64_KANAN) AND (i_pixel_row >G64_ATAS) AND (i_pixel_row < G64_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G65_KIRI) AND (i_pixel_column < G65_KANAN) AND (i_pixel_row > G65_ATAS) AND (i_pixel_row < G65_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G66_KIRI) AND (i_pixel_column < G66_KANAN) AND (i_pixel_row > G66_ATAS) AND (i_pixel_row < G66_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G67_KIRI) AND (i_pixel_column < G67_KANAN) AND (i_pixel_row > G67_ATAS) AND (i_pixel_row < G67_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G68_KIRI) AND (i_pixel_column < G68_KANAN) AND (i_pixel_row > G68_ATAS) AND (i_pixel_row < G68_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";		
		ELSIF ((i_pixel_column > G69_KIRI) AND (i_pixel_column < G69_KANAN) AND (i_pixel_row > G69_ATAS) AND (i_pixel_row < G69_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G70_KIRI) AND (i_pixel_column < G70_KANAN) AND (i_pixel_row > G70_ATAS) AND (i_pixel_row < G70_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G71_KIRI) AND (i_pixel_column < G71_KANAN) AND (i_pixel_row > G71_ATAS) AND (i_pixel_row < G71_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G72_KIRI) AND (i_pixel_column < G72_KANAN) AND (i_pixel_row > G72_ATAS) AND (i_pixel_row < G72_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G73_KIRI) AND (i_pixel_column < G73_KANAN) AND (i_pixel_row > G73_ATAS) AND (i_pixel_row < G73_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G74_KIRI) AND (i_pixel_column < G74_KANAN) AND (i_pixel_row > G74_ATAS) AND (i_pixel_row < G74_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G75_KIRI) AND (i_pixel_column < G75_KANAN) AND (i_pixel_row > G75_ATAS) AND (i_pixel_row < G75_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G76_KIRI) AND (i_pixel_column < G76_KANAN) AND (i_pixel_row > G76_ATAS) AND (i_pixel_row < G76_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G77_KIRI) AND (i_pixel_column < G77_KANAN) AND (i_pixel_row > G77_ATAS) AND (i_pixel_row < G77_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G78_KIRI) AND (i_pixel_column < G78_KANAN) AND (i_pixel_row > G78_ATAS) AND (i_pixel_row < G78_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G79_KIRI) AND (i_pixel_column < G79_KANAN) AND (i_pixel_row > G79_ATAS) AND (i_pixel_row < G79_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G80_KIRI) AND (i_pixel_column < G80_KANAN) AND (i_pixel_row > G80_ATAS) AND (i_pixel_row < G80_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G81_KIRI) AND (i_pixel_column < G81_KANAN) AND (i_pixel_row > G81_ATAS) AND (i_pixel_row < G81_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G82_KIRI) AND (i_pixel_column < G82_KANAN) AND (i_pixel_row > G82_ATAS) AND (i_pixel_row < G82_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G83_KIRI) AND (i_pixel_column < G83_KANAN) AND (i_pixel_row > G83_ATAS) AND (i_pixel_row < G83_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";		
		ELSIF ((i_pixel_column > G84_KIRI) AND (i_pixel_column < G84_KANAN) AND (i_pixel_row > G84_ATAS) AND (i_pixel_row < G84_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G85_KIRI) AND (i_pixel_column < G85_KANAN) AND (i_pixel_row > G85_ATAS) AND (i_pixel_row < G85_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G86_KIRI) AND (i_pixel_column < G86_KANAN) AND (i_pixel_row > G86_ATAS) AND (i_pixel_row < G86_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G87_KIRI) AND (i_pixel_column < G87_KANAN) AND (i_pixel_row > G87_ATAS) AND (i_pixel_row < G87_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G88_KIRI) AND (i_pixel_column < G88_KANAN) AND (i_pixel_row > G88_ATAS) AND (i_pixel_row < G88_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G89_KIRI) AND (i_pixel_column < G89_KANAN) AND (i_pixel_row > G89_ATAS) AND (i_pixel_row < G89_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G90_KIRI) AND (i_pixel_column < G90_KANAN) AND (i_pixel_row > G90_ATAS) AND (i_pixel_row < G90_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G91_KIRI) AND (i_pixel_column < G91_KANAN) AND (i_pixel_row > G91_ATAS) AND (i_pixel_row < G91_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G92_KIRI) AND (i_pixel_column < G92_KANAN) AND (i_pixel_row > G92_ATAS) AND (i_pixel_row < G92_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G93_KIRI) AND (i_pixel_column < G93_KANAN) AND (i_pixel_row > G93_ATAS) AND (i_pixel_row < G93_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G94_KIRI) AND (i_pixel_column < G94_KANAN) AND (i_pixel_row > G94_ATAS) AND (i_pixel_row < G94_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G95_KIRI) AND (i_pixel_column < G95_KANAN) AND (i_pixel_row > G95_ATAS) AND (i_pixel_row < G95_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G96_KIRI) AND (i_pixel_column < G96_KANAN) AND (i_pixel_row > G96_ATAS) AND (i_pixel_row < G96_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G97_KIRI) AND (i_pixel_column < G97_KANAN) AND (i_pixel_row > G97_ATAS) AND (i_pixel_row < G97_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G98_KIRI) AND (i_pixel_column < G98_KANAN) AND (i_pixel_row > G98_ATAS) AND (i_pixel_row < G98_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G99_KIRI) AND (i_pixel_column < G99_KANAN) AND (i_pixel_row > G99_ATAS) AND (i_pixel_row < G99_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G100_KIRI) AND (i_pixel_column < G100_KANAN) AND (i_pixel_row > G100_ATAS) AND (i_pixel_row < G100_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G101_KIRI) AND (i_pixel_column < G101_KANAN) AND (i_pixel_row > G101_ATAS) AND (i_pixel_row < G101_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G102_KIRI) AND (i_pixel_column < G102_KANAN) AND (i_pixel_row > G102_ATAS) AND (i_pixel_row < G102_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G103_KIRI) AND (i_pixel_column < G103_KANAN) AND (i_pixel_row > G103_ATAS) AND (i_pixel_row < G103_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G104_KIRI) AND (i_pixel_column < G104_KANAN) AND (i_pixel_row > G104_ATAS) AND (i_pixel_row < G104_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
			
		ELSE
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";
	END IF;
END IF;

--PENGAKTIFAN LAYAR UTAMA
IF i_K_BT = '0' AND (LEVEL = 1 OR LEVEL = 2) THEN
	UTAMA := TRUE;
END IF;

--LEVEL
IF i_K_BT = '1' AND LEVEL = 1 AND MENANG = FALSE AND KALAH1 = FALSE THEN --LEVEL 1

	IF clock40hz'event and clock40hz = '1' THEN
		KECEPATAN1 	:= 5;
		
	--WAKTU
	IF B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
		G62_ATAS	:= G62_ATAS;
		G62A_ATAS	:= G62A_ATAS;
		G62B_ATAS	:= G62B_ATAS;
		ELSE
			G62_ATAS	:= G62_ATAS + 1;
	IF G62_ATAS >= G62_BAWAH THEN
		G62_ATAS	:= G62_BAWAH;
		G62A_ATAS	:= G62A_ATAS + 1;
		END IF;
	IF G62A_ATAS >= G62A_BAWAH THEN
		G62A_ATAS	:= G62A_BAWAH;
		G62B_ATAS	:= G62B_ATAS + 1;
		END IF;
		END IF;
		
	--KONDISI KALAH
	IF G62B_ATAS >= G62B_BAWAH THEN
		G62B_ATAS 	:= G62B_ATAS;
		KALAH1		:= TRUE;
		END IF;
		
	--PAUSE
	IF i_K_BT = '0' AND LEVEL = 1 THEN
		KECEPATAN1 	:= 0;
		G62_ATAS	:= G62_ATAS;
		G62A_ATAS 	:= G62A_ATAS;
		G62B_ATAS 	:= G62B_ATAS;
		END IF;		
	
	--FINISH
	IF B1_KANAN <= F_KANAN AND B1_KIRI >= F_KIRI AND B1_ATAS >= F_ATAS AND B1_BAWAH <= F_BAWAH THEN
		LEVEL		:= 2;
		END IF;
	END IF;

	IF clock40hz'event and clock40hz = '1' AND i_M_US = '0' AND i_K_US = '1' AND i_H_US = '1' AND i_M_BT = '1' THEN
		B1_ATAS 	:= B1_ATAS - KECEPATAN1;   ---Arah Naik
		B1_BAWAH 	:= B1_BAWAH - KECEPATAN1;

		IF B1_ATAS <= 0 THEN
			B1_ATAS := 0;
			B1_BAWAH := 49;
			END IF;
		
		--GR2
		IF B1_ATAS <= GR2_BAWAH THEN
			B1_ATAS := GR2_BAWAH;
			B1_BAWAH := GR2_BAWAH + 50;
			END IF;
			
		--BATAS GC1
		IF B1_ATAS <= GC1_BAWAH AND B1_ATAS >= GC1_ATAS AND B1_KIRI < GC1_KANAN AND B1_KANAN > GC1_KIRI THEN
			B1_ATAS := GC1_BAWAH;
			B1_BAWAH := GC1_BAWAH + 50;
			END IF;

		--BATAS GC2
		IF B1_ATAS <= GC2_BAWAH AND B1_ATAS >= GC2_ATAS AND B1_KIRI < GC2_KANAN AND B1_KANAN > GC2_KIRI THEN
			B1_ATAS := GC2_BAWAH;
			B1_BAWAH := GC2_BAWAH + 50;
			END IF;
		
		--BATAS GC3
		IF B1_ATAS <= GC3_BAWAH AND B1_ATAS >= GC3_ATAS AND B1_KIRI < GC3_KANAN AND B1_KANAN > GC3_KIRI THEN
			B1_ATAS := GC3_BAWAH;
			B1_BAWAH := GC3_BAWAH + 50;
			END IF;
			
		--BATAS GC8
		IF B1_ATAS <= GC8_BAWAH AND B1_ATAS >= GC8_ATAS AND B1_KIRI < GC8_KANAN AND B1_KANAN > GC8_KIRI THEN
			B1_ATAS := GC8_BAWAH;
			B1_BAWAH := GC8_BAWAH + 50;
			END IF;
		
		--BATAS GC4
		IF B1_ATAS <= GC4_BAWAH AND B1_ATAS >= GC4_ATAS AND B1_KIRI < GC4_KANAN AND B1_KANAN > GC4_KIRI THEN
			B1_ATAS := GC4_BAWAH;
			B1_BAWAH := GC4_BAWAH + 50;
			END IF;
			
		--BATAS GR5
		IF B1_ATAS <= GR5_BAWAH AND B1_ATAS >= GR5_ATAS AND B1_KIRI < GR5_KANAN AND B1_KANAN > GR5_KIRI THEN
			B1_ATAS := GR5_BAWAH;
			B1_BAWAH := GR5_BAWAH + 50;
			END IF;
		
		--BATAS GR6
		IF B1_ATAS <= GR6_BAWAH AND B1_ATAS >= GR6_ATAS AND B1_KIRI < GR6_KANAN AND B1_KANAN > GR6_KIRI THEN

			B1_ATAS := GR6_BAWAH;
			B1_BAWAH := GR6_BAWAH + 50;
			END IF;
		
		--BATAS GR8
		IF B1_ATAS <= GR8_BAWAH AND B1_ATAS >= GR8_ATAS AND B1_KIRI < GR8_KANAN AND B1_KANAN > GR8_KIRI THEN
			B1_ATAS := GR8_BAWAH;
			B1_BAWAH := GR8_BAWAH + 50;
			END IF;
		
		--BATAS GR9
		IF B1_ATAS <= GR9_BAWAH AND B1_ATAS >= GR9_ATAS AND B1_KIRI < GR9_KANAN AND B1_KANAN > GR9_KIRI THEN
			B1_ATAS := GR9_BAWAH;
			B1_BAWAH := GR9_BAWAH + 50;
			END IF;
		
		
		--BATAS GR10
		IF B1_ATAS <= GR10_BAWAH AND B1_ATAS >= GR10_ATAS AND B1_KIRI < GR10_KANAN AND B1_KANAN > GR10_KIRI THEN
			B1_ATAS := GR10_BAWAH;
			B1_BAWAH := GR10_BAWAH + 50;
			END IF;
		
		--BATAS GR11
		IF B1_ATAS <= GR11_BAWAH AND B1_ATAS >= GR11_ATAS AND B1_KIRI < GR11_KANAN AND B1_KANAN > GR11_KIRI THEN
			B1_ATAS := GR11_BAWAH;
			B1_BAWAH := GR11_BAWAH + 50;
			END IF;
		
		--BATAS GR12
		IF B1_ATAS <= GR12_BAWAH AND B1_ATAS >= GR12_ATAS AND B1_KIRI < GR12_KANAN AND B1_KANAN > GR12_KIRI THEN
			B1_ATAS := GR12_BAWAH;
			B1_BAWAH := GR12_BAWAH + 50;
			END IF;
			
		--BATAS GR13
		IF B1_ATAS <= GR13_BAWAH AND B1_ATAS >= GR13_ATAS AND B1_KIRI < GR13_KANAN AND B1_KANAN > GR13_KIRI THEN
			B1_ATAS := GR13_BAWAH;
			B1_BAWAH := GR13_BAWAH + 50;
			END IF;
		
		--BATAS GR14
		IF B1_ATAS <= GR14_BAWAH AND B1_ATAS >= GR14_ATAS AND B1_KIRI < GR14_KANAN AND B1_KANAN > GR14_KIRI THEN
			B1_ATAS := GR14_BAWAH;
			B1_BAWAH := GR14_BAWAH + 50;
			END IF;
			
	ELSIF clock40hz'event and clock40hz = '1' AND i_M_US = '1' AND i_K_US = '0' AND i_H_US = '1' AND i_M_BT = '1' THEN
		B1_ATAS 	:= B1_ATAS + KECEPATAN1;    ---Arah Turun
		B1_BAWAH	:= B1_BAWAH + KECEPATAN1;
		
		IF B1_BAWAH >= 479 THEN
			B1_ATAS := 479 -49;
			B1_BAWAH := 479;
			END IF;
		
		--GR3
		IF B1_BAWAH >= GR3_ATAS THEN
			B1_ATAS := GR3_ATAS - 50;
			B1_BAWAH := GR3_ATAS;
			END IF;
			
		--BATAS GC8
		IF B1_BAWAH >= GC8_ATAS AND B1_BAWAH <= GC8_BAWAH AND B1_KIRI < GC8_KANAN AND B1_KANAN > GC8_KIRI THEN
			B1_ATAS := GC8_ATAS - 50;
			B1_BAWAH := GC8_ATAS;
			END IF;

		--BATAS GC5
		IF B1_BAWAH >= GC5_ATAS AND B1_BAWAH <= GC5_BAWAH AND B1_KIRI < GC5_KANAN AND B1_KANAN > GC5_KIRI THEN
			B1_ATAS := GC5_ATAS - 50;
			B1_BAWAH := GC5_ATAS;
			END IF;

		--BATAS GC4
		IF B1_BAWAH >= GC4_ATAS AND B1_BAWAH <= GC4_BAWAH AND B1_KIRI < GC4_KANAN AND B1_KANAN > GC4_KIRI THEN
			B1_ATAS := GC4_ATAS - 50;
			B1_BAWAH := GC4_ATAS;
			END IF;

		--BATAS GC7
		IF B1_BAWAH >= GC7_ATAS AND B1_BAWAH <= GC7_BAWAH AND B1_KIRI < GC7_KANAN AND B1_KANAN > GC7_KIRI THEN
			B1_ATAS := GC7_ATAS - 50;
			B1_BAWAH := GC7_ATAS;
			END IF;
			
		--BATAS GC8
		IF B1_BAWAH >= GC8_ATAS AND B1_BAWAH <= GC8_BAWAH AND B1_KIRI < GC8_KANAN AND B1_KANAN > GC8_KIRI THEN
			B1_ATAS := GC8_ATAS - 50;
			B1_BAWAH := GC8_ATAS;
			END IF;
			
						
		--BATAS GR5
		IF B1_BAWAH >= GR5_ATAS AND B1_BAWAH <= GR5_BAWAH AND B1_KIRI < GR5_KANAN AND B1_KANAN > GR5_KIRI THEN
			B1_ATAS := GR5_ATAS - 50;
			B1_BAWAH := GR5_ATAS;
			END IF;
			
		--BATAS GR6
		IF B1_BAWAH >= GR6_ATAS AND B1_BAWAH <= GR6_BAWAH AND B1_KIRI < GR6_KANAN AND B1_KANAN > GR6_KIRI THEN
			B1_ATAS := GR6_ATAS - 50;
			B1_BAWAH := GR6_ATAS;
			END IF;


		--BATAS GR8
		IF B1_BAWAH >= GR8_ATAS AND B1_BAWAH <= GR8_BAWAH AND B1_KIRI < GR8_KANAN AND B1_KANAN > GR8_KIRI THEN
			B1_ATAS := GR8_ATAS - 50;
			B1_BAWAH := GR8_ATAS;
			END IF;

		--BATAS GR9
		IF B1_BAWAH >= GR9_ATAS AND B1_BAWAH <= GR9_BAWAH AND B1_KIRI < GR9_KANAN AND B1_KANAN > GR9_KIRI THEN
			B1_ATAS := GR9_ATAS - 50;
			B1_BAWAH := GR9_ATAS;
			END IF;
			
		--BATAS GR10
		IF B1_BAWAH >= GR10_ATAS AND B1_BAWAH <= GR10_BAWAH AND B1_KIRI < GR10_KANAN AND B1_KANAN > GR10_KIRI THEN
			B1_ATAS := GR10_ATAS - 50;
			B1_BAWAH := GR10_ATAS;
			END IF;
		
		--BATAS GR11
		IF B1_BAWAH >= GR11_ATAS AND B1_BAWAH <= GR11_BAWAH AND B1_KIRI < GR11_KANAN AND B1_KANAN > GR11_KIRI THEN
			B1_ATAS := GR11_ATAS - 50;
			B1_BAWAH := GR11_ATAS;
			END IF;
			
		--BATAS GR14
		IF B1_BAWAH >= GR14_ATAS AND B1_BAWAH <= GR14_BAWAH AND B1_KIRI < GR14_KANAN AND B1_KANAN > GR14_KIRI THEN
			B1_ATAS := GR14_ATAS - 50;
			B1_BAWAH := GR14_ATAS;
			END IF;

	ELSIF clock40hz'event and clock40hz = '1' AND i_M_US = '1' AND i_K_US = '1' AND i_H_US = '0' AND i_M_BT = '1' THEN
		B1_KANAN 	:= B1_KANAN + KECEPATAN1;  ---Arah kanan
		B1_KIRI 	:= B1_KIRI + KECEPATAN1;
		
		IF B1_KANAN >= 639 THEN
			B1_KANAN := 639;
			B1_KIRI := 639 -49;
			END IF;
			
		--GR4
		IF B1_KANAN >= GR4_KIRI THEN
			B1_KIRI := GR4_KIRI - 50;
			B1_KANAN := GR4_KIRI;
			END IF;
		
		--BATAS GC1
		IF B1_KANAN >= GC1_KIRI AND B1_KANAN <= GC1_KANAN AND B1_BAWAH > GC1_ATAS AND B1_ATAS < GC1_BAWAH THEN
			B1_KANAN := GC1_KIRI;
			B1_KIRI := GC1_KIRI - 50;
			END IF;
		
		--BATAS GC2
		IF B1_KANAN >= GC2_KIRI AND B1_KANAN <= GC2_KANAN AND B1_BAWAH > GC2_ATAS AND B1_ATAS < GC2_BAWAH THEN
			B1_KANAN := GC2_KIRI;
			B1_KIRI := GC2_KIRI - 50;
			END IF;
			
		--BATAS GC3
		IF B1_KANAN >= GC3_KIRI AND B1_KANAN <= GC3_KANAN AND B1_BAWAH > GC3_ATAS AND B1_ATAS < GC3_BAWAH THEN
			B1_KANAN := GC3_KIRI;
			B1_KIRI := GC3_KIRI - 50;
			END IF;
			
		--BATAS GC8
		IF B1_KANAN >= GC8_KIRI AND B1_KANAN <= GC8_KANAN AND B1_BAWAH > GC8_ATAS AND B1_ATAS < GC8_BAWAH THEN
			B1_KANAN := GC8_KIRI;
			B1_KIRI := GC8_KIRI - 50;
			END IF;
		
		--BATAS GC4
		IF B1_KANAN >= GC4_KIRI AND B1_KANAN <= GC4_KANAN AND B1_BAWAH > GC4_ATAS AND B1_ATAS < GC4_BAWAH THEN
			B1_KANAN := GC4_KIRI;
			B1_KIRI := GC4_KIRI - 50;
			END IF;
			
		--BATAS GC5
		IF B1_KANAN >= GC5_KIRI AND B1_KANAN <= GC5_KANAN AND B1_BAWAH > GC5_ATAS AND B1_ATAS < GC5_BAWAH THEN
			B1_KANAN := GC5_KIRI;
			B1_KIRI := GC5_KIRI - 50;
			END IF;
		
		--BATAS GC7
		IF B1_KANAN >= GC7_KIRI AND B1_KANAN <= GC7_KANAN AND B1_BAWAH > GC7_ATAS AND B1_ATAS < GC7_BAWAH THEN
			B1_KANAN := GC7_KIRI;
			B1_KIRI := GC7_KIRI - 50;
			END IF;
			
		--BATAS GR9
		IF B1_KANAN >= GR9_KIRI AND B1_KANAN <= GR9_KANAN AND B1_BAWAH > GR9_ATAS AND B1_ATAS < GR9_BAWAH THEN
			B1_KANAN := GR9_KIRI;
			B1_KIRI := GR9_KIRI - 50;
			END IF;
		
		--BATAS GR10
		IF B1_KANAN >= GR10_KIRI AND B1_KANAN <= GR10_KANAN AND B1_BAWAH > GR10_ATAS AND B1_ATAS < GR10_BAWAH THEN
			B1_KANAN := GR10_KIRI;
			B1_KIRI := GR10_KIRI - 50;
			END IF;
		
		--BATAS GR14
		IF B1_KANAN >= GR14_KIRI AND B1_KANAN <= GR14_KANAN AND B1_BAWAH > GR14_ATAS AND B1_ATAS < GR14_BAWAH THEN
			B1_KANAN := GR14_KIRI;
			B1_KIRI := GR14_KIRI - 50;
			END IF;		

	ELSIF clock40hz'event and clock40hz = '1' AND i_M_US = '1' AND i_K_US = '1' AND i_H_US = '1' AND i_M_BT = '0' THEN
		B1_KANAN 	:= B1_KANAN - KECEPATAN1;  ---Arah Kiri
		B1_KIRI 	:= B1_KIRI - KECEPATAN1;
		
		IF B1_KIRI <= 0 THEN
			B1_KIRI := 0;
			B1_KANAN := 49;
			END IF;	
	
		--GR1
		IF B1_KIRI <= GR1_KANAN THEN
			B1_KIRI := GR1_KANAN;
			B1_KANAN := GR1_KANAN + 50;
			END IF;
	
		--BATAS GC1
		IF B1_KIRI <= GC1_KANAN AND B1_KIRI >= GC1_KIRI AND B1_ATAS < GC1_BAWAH  AND B1_BAWAH > GC1_ATAS THEN
			B1_KIRI := GC1_KANAN;
			B1_KANAN := GC1_KANAN + 50;
			END IF;
	
		--BATAS GC2
		IF B1_KIRI <= GC2_KANAN AND B1_KIRI >= GC2_KIRI AND B1_ATAS < GC2_BAWAH  AND B1_BAWAH > GC2_ATAS THEN
			B1_KIRI := GC2_KANAN;
			B1_KANAN := GC2_KANAN + 50;
			END IF;
	
		--BATAS GC3
		IF B1_KIRI <= GC3_KANAN AND B1_KIRI >= GC3_KIRI AND B1_ATAS < GC3_BAWAH  AND B1_BAWAH > GC3_ATAS THEN
			B1_KIRI := GC3_KANAN;
			B1_KANAN := GC3_KANAN + 50;
			END IF;
			
		--BATAS GC8
		IF B1_KIRI <= GC8_KANAN AND B1_KIRI >= GC8_KIRI AND B1_ATAS < GC8_BAWAH  AND B1_BAWAH > GC8_ATAS THEN
			B1_KIRI := GC8_KANAN;
			B1_KANAN := GC8_KANAN + 50;
			END IF;
	
	
		--BATAS GC4
		IF B1_KIRI <= GC4_KANAN AND B1_KIRI >= GC4_KIRI AND B1_ATAS < GC4_BAWAH  AND B1_BAWAH > GC4_ATAS THEN
			B1_KIRI := GC4_KANAN;
			B1_KANAN := GC4_KANAN + 50;
			END IF;
	
		--BATAS GC5
		IF B1_KIRI <= GC5_KANAN AND B1_KIRI >= GC5_KIRI AND B1_ATAS < GC5_BAWAH  AND B1_BAWAH > GC5_ATAS THEN
			B1_KIRI := GC5_KANAN;
			B1_KANAN := GC5_KANAN + 50;
			END IF;
	
		--BATAS GC7
		IF B1_KIRI <= GC7_KANAN AND B1_KIRI >= GC7_KIRI AND B1_ATAS < GC7_BAWAH  AND B1_BAWAH > GC7_ATAS THEN
			B1_KIRI := GC7_KANAN;
			B1_KANAN := GC7_KANAN + 50;
			END IF;
	
		--BATAS GR5
		IF B1_KIRI <= GR5_KANAN AND B1_KIRI >= GR5_KIRI AND B1_ATAS < GR5_BAWAH  AND B1_BAWAH > GR5_ATAS THEN
			B1_KIRI := GR5_KANAN;
			B1_KANAN := GR5_KANAN + 50;
			END IF;
	
		--BATAS GR6
		IF B1_KIRI <= GR6_KANAN AND B1_KIRI >= GR6_KIRI AND B1_ATAS < GR6_BAWAH  AND B1_BAWAH > GR6_ATAS THEN
			B1_KIRI := GR6_KANAN;
			B1_KANAN := GR6_KANAN + 50;
			END IF;
			
		--BATAS GR8
		IF B1_KIRI <= GR8_KANAN AND B1_KIRI >= GR8_KIRI AND B1_ATAS < GR8_BAWAH  AND B1_BAWAH > GR8_ATAS THEN
			B1_KIRI := GR8_KANAN;
			B1_KANAN := GR8_KANAN + 50;
			END IF;
			
		--BATAS GR9
		IF B1_KIRI <= GR9_KANAN AND B1_KIRI >= GR9_KIRI AND B1_ATAS < GR9_BAWAH  AND B1_BAWAH > GR9_ATAS THEN
			B1_KIRI := GR9_KANAN;
			B1_KANAN := GR9_KANAN + 50;
			END IF;
			
		--BATAS GR10
		IF B1_KIRI <= GR10_KANAN AND B1_KIRI >= GR10_KIRI AND B1_ATAS < GR10_BAWAH  AND B1_BAWAH > GR10_ATAS THEN
			B1_KIRI := GR10_KANAN;
			B1_KANAN := GR10_KANAN + 50;
			END IF;
			
		--BATAS GR11
		IF B1_KIRI <= GR11_KANAN AND B1_KIRI >= GR11_KIRI AND B1_ATAS < GR11_BAWAH  AND B1_BAWAH > GR11_ATAS THEN
			B1_KIRI := GR11_KANAN;
			B1_KANAN := GR11_KANAN + 50;
			END IF;
		--BATAS GR12
		IF B1_KIRI <= GR12_KANAN AND B1_KIRI >= GR12_KIRI AND B1_ATAS < GR12_BAWAH  AND B1_BAWAH > GR12_ATAS THEN
			B1_KIRI := GR12_KANAN;
			B1_KANAN := GR12_KANAN + 50;
			END IF;
		--BATAS GR13
		IF B1_KIRI <= GR13_KANAN AND B1_KIRI >= GR13_KIRI AND B1_ATAS < GR13_BAWAH  AND B1_BAWAH > GR13_ATAS THEN
			B1_KIRI := GR13_KANAN;
			B1_KANAN := GR13_KANAN + 50;
			END IF;
		--BATAS GR14
		IF B1_KIRI <= GR14_KANAN AND B1_KIRI >= GR14_KIRI AND B1_ATAS < GR14_BAWAH  AND B1_BAWAH > GR14_ATAS THEN
			B1_KIRI := GR14_KANAN;
			B1_KANAN := GR14_KANAN + 50;
			END IF;
	
ELSE

B1_KIRI := B1_KIRI;
B1_KANAN := B1_KANAN;
B1_BAWAH := B1_BAWAH;
B1_ATAS := B1_ATAS;


END IF;


IF ((i_pixel_column > B1_KIRI) AND (i_pixel_column < B1_KANAN) AND (i_pixel_row >B1_ATAS) AND (i_pixel_row < B1_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"00"; o_blue <= X"00";
						
		ELSIF ((i_pixel_column > GR1_KIRI) AND (i_pixel_column < GR1_KANAN) AND (i_pixel_row > GR1_ATAS) AND (i_pixel_row < GR1_BAWAH)) THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GR2_KIRI) AND (i_pixel_column < GR2_KANAN) AND (i_pixel_row > GR2_ATAS) AND (i_pixel_row < GR2_BAWAH)) THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GR3_KIRI) AND (i_pixel_column < GR3_KANAN) AND (i_pixel_row > GR3_ATAS) AND (i_pixel_row < GR3_BAWAH)) THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GR4_KIRI) AND (i_pixel_column < GR4_KANAN) AND (i_pixel_row > GR4_ATAS) AND (i_pixel_row < GR4_BAWAH)) THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GR5_KIRI) AND (i_pixel_column < GR5_KANAN) AND (i_pixel_row > GR5_ATAS) AND (i_pixel_row < GR5_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GR6_KIRI) AND (i_pixel_column < GR6_KANAN) AND (i_pixel_row > GR6_ATAS) AND (i_pixel_row < GR6_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GR8_KIRI) AND (i_pixel_column < GR8_KANAN) AND (i_pixel_row > GR8_ATAS) AND (i_pixel_row < GR8_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";
		ELSIF ((i_pixel_column > GR9_KIRI) AND (i_pixel_column < GR9_KANAN) AND (i_pixel_row > GR9_ATAS) AND (i_pixel_row < GR9_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GR10_KIRI) AND (i_pixel_column < GR10_KANAN) AND (i_pixel_row > GR10_ATAS) AND (i_pixel_row < GR10_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GR11_KIRI) AND (i_pixel_column < GR11_KANAN) AND (i_pixel_row > GR11_ATAS) AND (i_pixel_row < GR11_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GR12_KIRI) AND (i_pixel_column < GR12_KANAN) AND (i_pixel_row > GR12_ATAS) AND (i_pixel_row < GR12_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GR13_KIRI) AND (i_pixel_column < GR13_KANAN) AND (i_pixel_row > GR13_ATAS) AND (i_pixel_row < GR13_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GR14_KIRI) AND (i_pixel_column < GR14_KANAN) AND (i_pixel_row > GR14_ATAS) AND (i_pixel_row < GR14_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";		
		ELSIF ((i_pixel_column > GC1_KIRI) AND (i_pixel_column < GC1_KANAN) AND (i_pixel_row > GC1_ATAS) AND (i_pixel_row < GC1_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";		
		ELSIF ((i_pixel_column > GC2_KIRI) AND (i_pixel_column < GC2_KANAN) AND (i_pixel_row > GC2_ATAS) AND (i_pixel_row < GC2_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GC3_KIRI) AND (i_pixel_column < GC3_KANAN) AND (i_pixel_row > GC3_ATAS) AND (i_pixel_row < GC3_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GC4_KIRI) AND (i_pixel_column < GC4_KANAN) AND (i_pixel_row > GC4_ATAS) AND (i_pixel_row < GC4_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GC5_KIRI) AND (i_pixel_column < GC5_KANAN) AND (i_pixel_row > GC5_ATAS) AND (i_pixel_row < GC5_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GC7_KIRI) AND (i_pixel_column < GC7_KANAN) AND (i_pixel_row > GC7_ATAS) AND (i_pixel_row < GC7_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > GC8_KIRI) AND (i_pixel_column < GC8_KANAN) AND (i_pixel_row > GC8_ATAS) AND (i_pixel_row < GC8_BAWAH)) AND B1_ATAS >= S_ATAS AND B1_KIRI >= S_KIRI AND B1_KANAN <= S_KANAN AND B1_BAWAH <= S_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";		
		ELSIF ((i_pixel_column > F_KIRI) AND (i_pixel_column < F_KANAN) AND (i_pixel_row > F_ATAS) AND (i_pixel_row < F_BAWAH)) THEN
			o_red <= X"64"; o_green <= X"FA"; o_blue <= X"C8";	
		
		--PERUBAHAN WARNA BATAS LEVEL 1	
		ELSIF ((i_pixel_column > GR5_KIRI) AND (i_pixel_column < GR5_KANAN) AND (i_pixel_row > GR5_ATAS) AND (i_pixel_row < GR5_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > GR6_KIRI) AND (i_pixel_column < GR6_KANAN) AND (i_pixel_row > GR6_ATAS) AND (i_pixel_row < GR6_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > GR8_KIRI) AND (i_pixel_column < GR8_KANAN) AND (i_pixel_row > GR8_ATAS) AND (i_pixel_row < GR8_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > GR9_KIRI) AND (i_pixel_column < GR9_KANAN) AND (i_pixel_row > GR9_ATAS) AND (i_pixel_row < GR9_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > GR10_KIRI) AND (i_pixel_column < GR10_KANAN) AND (i_pixel_row > GR10_ATAS) AND (i_pixel_row < GR10_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > GR11_KIRI) AND (i_pixel_column < GR11_KANAN) AND (i_pixel_row > GR11_ATAS) AND (i_pixel_row < GR11_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > GR12_KIRI) AND (i_pixel_column < GR12_KANAN) AND (i_pixel_row > GR12_ATAS) AND (i_pixel_row < GR12_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > GR13_KIRI) AND (i_pixel_column < GR13_KANAN) AND (i_pixel_row > GR13_ATAS) AND (i_pixel_row < GR13_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > GR14_KIRI) AND (i_pixel_column < GR14_KANAN) AND (i_pixel_row > GR14_ATAS) AND (i_pixel_row < GR14_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";		
		ELSIF ((i_pixel_column > GC1_KIRI) AND (i_pixel_column < GC1_KANAN) AND (i_pixel_row > GC1_ATAS) AND (i_pixel_row < GC1_BAWAH))  THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";		
		ELSIF ((i_pixel_column > GC2_KIRI) AND (i_pixel_column < GC2_KANAN) AND (i_pixel_row > GC2_ATAS) AND (i_pixel_row < GC2_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > GC3_KIRI) AND (i_pixel_column < GC3_KANAN) AND (i_pixel_row > GC3_ATAS) AND (i_pixel_row < GC3_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > GC4_KIRI) AND (i_pixel_column < GC4_KANAN) AND (i_pixel_row > GC4_ATAS) AND (i_pixel_row < GC4_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > GC5_KIRI) AND (i_pixel_column < GC5_KANAN) AND (i_pixel_row > GC5_ATAS) AND (i_pixel_row < GC5_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > GC7_KIRI) AND (i_pixel_column < GC7_KANAN) AND (i_pixel_row > GC7_ATAS) AND (i_pixel_row < GC7_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > GC8_KIRI) AND (i_pixel_column < GC8_KANAN) AND (i_pixel_row > GC8_ATAS) AND (i_pixel_row < GC8_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
			
		--WAKTU
		ELSIF ((i_pixel_column > G62_KIRI) AND (i_pixel_column < G62_KANAN) AND (i_pixel_row > G62_ATAS) AND (i_pixel_row < G62_BAWAH)) THEN
			o_red <= X"00"; o_green <= X"FF"; o_blue <= X"00";
		ELSIF ((i_pixel_column > G62A_KIRI) AND (i_pixel_column < G62A_KANAN) AND (i_pixel_row > G62A_ATAS) AND (i_pixel_row < G62A_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"00";
		ELSIF ((i_pixel_column > G62B_KIRI) AND (i_pixel_column < G62B_KANAN) AND (i_pixel_row > G62B_ATAS) AND (i_pixel_row < G62B_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"00"; o_blue <= X"00";
			
		ELSE 
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
	END IF;

ELSIF i_K_BT = '1' AND LEVEL = 2 AND MENANG = FALSE AND KALAH = FALSE THEN --LEVEL 2

	IF clock40hz'event and clock40hz = '1' THEN
		KECEPATAN	:= 5;
		
	--WAKTU
	IF B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
		G63_ATAS	:= G63_ATAS;
		G63A_ATAS	:= G63A_ATAS;
		G63B_ATAS	:= G63B_ATAS;
		ELSE
			G63_ATAS	:= G63_ATAS + 1;
	IF G63_ATAS >= G63_BAWAH THEN
		G63_ATAS 	:= G63_BAWAH;
		G63A_ATAS	:= G63A_ATAS + 1;
		END IF;
	IF G63A_ATAS >= G63A_BAWAH THEN
		G63A_ATAS	:= G63A_BAWAH;
		G63B_ATAS 	:= G63B_ATAS + 1;
		END IF;
		END IF;
			
	--KONDISI KALAH
	IF G63B_ATAS >= G63B_BAWAH THEN
		G63B_ATAS 	:= G63B_ATAS;
		KALAH		:= TRUE;
		END IF;
		
	--PAUSE
	IF i_K_BT = '0' AND LEVEL = 2 THEN
		KECEPATAN 	:= 0;
		G63_ATAS 	:= G63_ATAS;
		G63A_ATAS 	:= G63A_ATAS;
		G63B_ATAS 	:= G63B_ATAS;
		END IF;
		
	--KONDISI MENANG
	IF B_KANAN <= G61_KANAN AND B_KIRI >= G61_KIRI AND B_ATAS >= G61_ATAS AND B_BAWAH <= G61_BAWAH THEN
		MENANG		:= TRUE;
		END IF;
	END IF;
	
	IF clock40hz'event and clock40hz = '1' AND i_M_US = '0' AND i_K_US = '1' AND i_H_US = '1' AND i_M_BT = '1' THEN
		B_ATAS 		:= B_ATAS - KECEPATAN;   ---Arah Naik
		B_BAWAH		:= B_BAWAH - KECEPATAN;

		IF B_ATAS <= 0 THEN
			B_ATAS := 0;
			B_BAWAH := 49;
			END IF;
		
	--BINGKAI ATAS
		IF B_ATAS <= G1_BAWAH THEN
			B_ATAS := G1_BAWAH;
			B_BAWAH := G1_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL I DAN M POJOK KIRI BAWAH
		IF B_ATAS <= G6_BAWAH AND B_ATAS >= G6_ATAS AND B_KIRI < G6_KANAN THEN
			B_ATAS := G6_BAWAH;
			B_BAWAH := G6_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL DI BAWAH M
		IF B_ATAS <= G13_BAWAH AND B_ATAS >= G13_ATAS AND B_KANAN > G13_KIRI AND B_KIRI < G13_KANAN  THEN
			B_ATAS := G13_BAWAH;
			B_BAWAH := G13_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL M DI POJOK KANAN BAWAH AMPE A
		IF B_ATAS <= G14_BAWAH AND B_ATAS >= G14_ATAS AND B_KANAN > G14_KIRI AND B_KIRI < G14_KANAN  THEN
			B_ATAS := G14_BAWAH;
			B_BAWAH := G14_BAWAH + 30;
			END IF;
	--KOTAK DI TENGAH A
		IF B_ATAS <= G16_BAWAH AND B_ATAS >= G16_ATAS AND B_KANAN > G16_KIRI AND B_KIRI < G16_KANAN  THEN
			B_ATAS := G16_BAWAH;
			B_BAWAH := G16_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL DI TENGAH A
		IF B_ATAS <= G17_BAWAH AND B_ATAS >= G17_ATAS AND B_KANAN > G17_KIRI AND B_KIRI < G17_KANAN  THEN
			B_ATAS := G17_BAWAH;
			B_BAWAH := G17_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL A DI POJOK KANAN BAWAH
		IF B_ATAS <= G18_BAWAH AND B_ATAS >= G18_ATAS AND B_KANAN > G18_KIRI AND B_KIRI < G18_KANAN  THEN
			B_ATAS := G18_BAWAH;
			B_BAWAH := G18_BAWAH + 30;
			END IF;
	--KOTAK DI BAWAH I
		IF B_ATAS <= G22_BAWAH AND B_ATAS >= G22_ATAS AND B_KANAN > G22_KIRI AND B_KIRI < G22_KANAN  THEN
			B_ATAS := G22_BAWAH;
			B_BAWAH := G22_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL_1 DI BAWAH I
		IF B_ATAS <= G23_BAWAH AND B_ATAS >= G23_ATAS AND B_KIRI < G23_KANAN  THEN
			B_ATAS := G23_BAWAH;
			B_BAWAH := G23_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL_2 DI BAWAH I
		IF B_ATAS <= G24_BAWAH AND B_ATAS >= G24_ATAS AND B_ATAS >= G24_ATAS AND B_KIRI < G24_KANAN  THEN
			B_ATAS := G24_BAWAH;
			B_BAWAH := G24_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL_3 DI BAWAH I
		IF B_ATAS <= G25_BAWAH AND B_ATAS >= G25_ATAS AND B_ATAS >= G25_ATAS AND B_KIRI < G25_KANAN  THEN
			B_ATAS := G25_BAWAH;
			B_BAWAH := G25_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL_1 DI BAWAH M
		IF B_ATAS <= G26_BAWAH AND B_ATAS >= G26_ATAS AND B_ATAS >= G26_ATAS AND B_KANAN > G26_KIRI AND B_KIRI < G26_KANAN  THEN
			B_ATAS := G26_BAWAH;
			B_BAWAH := G26_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL_2 DI BAWAH M
		IF B_ATAS <= G30_BAWAH AND B_ATAS >= G30_ATAS AND B_ATAS >= G30_ATAS AND B_KANAN > G30_KIRI AND B_KIRI < G30_KANAN  THEN
			B_ATAS := G30_BAWAH;
			B_BAWAH := G30_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL_3 DI BAWAH M
		IF B_ATAS <= G31_BAWAH AND B_ATAS >= G31_ATAS AND B_KANAN > G31_KIRI AND B_KIRI < G31_KANAN  THEN
			B_ATAS := G31_BAWAH;
			B_BAWAH := G31_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL DI BAWAH A
		IF B_ATAS <= G32_BAWAH AND B_ATAS >= G32_ATAS AND B_KANAN > G32_KIRI AND B_KIRI < G32_KANAN  THEN
			B_ATAS := G32_BAWAH;
			B_BAWAH := G32_BAWAH + 30;
			END IF;
	--KOTAK DI BAWAH A
		IF B_ATAS <= G33_BAWAH AND B_ATAS >= G33_ATAS AND B_KANAN > G33_KIRI AND B_KIRI < G33_KANAN  THEN
			B_ATAS := G33_BAWAH;
			B_BAWAH := G33_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL DI KANAN A
		IF B_ATAS <= G37_BAWAH AND B_ATAS >= G37_ATAS AND B_KANAN > G37_KIRI AND B_KIRI < G37_KANAN  THEN
			B_ATAS := G37_BAWAH;
			B_BAWAH := G37_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL_1 DI BAWAH U
		IF B_ATAS <= G42_BAWAH AND B_ATAS >= G42_ATAS AND B_KANAN > G42_KIRI AND B_KIRI < G42_KANAN  THEN
			B_ATAS := G42_BAWAH;
			B_BAWAH := G42_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL_3 DI BAWAH U
		IF B_ATAS <= G44_BAWAH AND B_ATAS >= G44_ATAS AND B_KANAN > G44_KIRI AND B_KIRI < G44_KANAN  THEN
			B_ATAS := G44_BAWAH;
			B_BAWAH := G44_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL_4 DI BAWAH U
		IF B_ATAS <= G45_BAWAH AND B_ATAS >= G45_ATAS AND B_KANAN > G45_KIRI AND B_KIRI < G45_KANAN  THEN
			B_ATAS := G45_BAWAH;
			B_BAWAH := G45_BAWAH + 30;
			END IF;
	--GARIS HORIZONTAL_5 DI BAWAH U
		IF B_ATAS <= G46_BAWAH AND B_ATAS >= G46_ATAS AND B_KANAN > G46_KIRI AND B_KIRI < G46_KANAN  THEN
			B_ATAS := G46_BAWAH;
			B_BAWAH := G46_BAWAH + 30;
			END IF;
	--TELEPORT 3
		IF B_KANAN <= G49_KANAN AND B_KIRI >= G49_KIRI AND B_ATAS >= G49_ATAS AND B_BAWAH <= G49_BAWAH THEN
			B_ATAS := 380;
			B_BAWAH := 380 + 30;
			B_KIRI := 10;
			B_KANAN := 10 + 30;
			END IF;
	--TELEPORT 12
		IF B_KANAN <= G58_KANAN AND B_KIRI >= G58_KIRI AND B_ATAS >= G58_ATAS AND B_BAWAH <= G58_BAWAH THEN
			B_ATAS := 130;
			B_BAWAH := 130 + 30;
			B_KIRI := 160;
			B_KANAN := 160 + 30;
			END IF;
	--TELEPORT 14
		IF B_KANAN <= G60_KANAN AND B_KIRI >= G60_KIRI AND B_ATAS >= G60_ATAS AND B_BAWAH <= G60_BAWAH THEN
			B_ATAS := 170;
			B_BAWAH := 170 + 30;
			B_KIRI := 10;
			B_KANAN := 10 + 30;
			END IF;
		
	ELSIF clock40hz'event and clock40hz = '1' AND i_M_US = '1' AND i_K_US = '0' AND i_H_US = '1' AND i_M_BT = '1' THEN
		B_ATAS 		:= B_ATAS + KECEPATAN;    ---Arah Turun
		B_BAWAH 	:= B_BAWAH + KECEPATAN;
		
		IF B_BAWAH >= 479 THEN
			B_ATAS := 479 -49;
			B_BAWAH := 479;
			END IF;
			
	--BINGKAI BAWAH
		IF B_BAWAH >= G3_ATAS THEN
			B_ATAS := G3_ATAS - 30;
			B_BAWAH := G3_ATAS;
			END IF;
	--GARIS HORIZONTAL DI ATAS KIRI M
		IF B_BAWAH >= G11_ATAS AND B_BAWAH <= G11_BAWAH AND B_KIRI < G11_KANAN AND B_KANAN > G11_KIRI THEN
			B_ATAS := G11_ATAS - 30;
			B_BAWAH := G11_ATAS;
			END IF;
	--GARIS HORIZONTAL DI ATAS KANAN M
		IF B_BAWAH >= G12_ATAS AND B_BAWAH <= G12_BAWAH AND B_KIRI < G12_KANAN AND B_KANAN > G12_KIRI THEN
			B_ATAS := G12_ATAS - 30;
			B_BAWAH := G12_ATAS;
			END IF;
	--GARIS HORIZONTAL M BAWAH
		IF B_BAWAH >= G13_ATAS AND B_BAWAH <= G13_BAWAH AND B_KIRI < G13_KANAN AND B_KANAN > G13_KIRI THEN
			B_ATAS := G13_ATAS - 30;
			B_BAWAH := G13_ATAS;
			END IF;
	--KOTAK DI TENGAH A
		IF B_BAWAH >= G16_ATAS AND B_BAWAH <= G16_BAWAH AND B_KIRI < G16_KANAN AND B_KANAN > G16_KIRI THEN
			B_ATAS := G16_ATAS - 30;
			B_BAWAH := G16_ATAS;
			END IF;
	--GARIS HORIZONTAL DI TENGAH A
		IF B_BAWAH >= G17_ATAS AND B_BAWAH <= G17_BAWAH AND B_KIRI < G17_KANAN AND B_KANAN > G17_KIRI THEN
			B_ATAS := G17_ATAS - 30;
			B_BAWAH := G17_ATAS;
			END IF;
	--GARIS HORIZONTAL_1 DI BAWAH I
		IF B_BAWAH >= G23_ATAS AND B_BAWAH <= G23_BAWAH AND B_KIRI < G23_KANAN THEN
			B_ATAS := G23_ATAS - 30;
			B_BAWAH := G23_ATAS;
			END IF;
	--GARIS HORIZONTAL_2 DI BAWAH I
		IF B_BAWAH >= G24_ATAS AND B_BAWAH <= G24_BAWAH AND B_KIRI < G24_KANAN THEN
			B_ATAS := G24_ATAS -30;
			B_BAWAH := G24_ATAS;
			END IF;
	--GARIS HORIZONTAL_3 DI BAWAH I
		IF B_BAWAH >= G25_ATAS AND B_BAWAH <= G25_BAWAH AND B_KIRI < G25_KANAN THEN
			B_ATAS := G25_ATAS - 30;
			B_BAWAH := G25_ATAS;
			END IF;
	--GARIS HORIZONTAL_1 DI BAWAH M
		IF B_BAWAH >= G26_ATAS AND B_BAWAH <= G26_BAWAH AND B_KIRI < G26_KANAN AND B_KANAN > G26_KIRI THEN
			B_ATAS := G26_ATAS - 30;
			B_BAWAH := G26_ATAS;
			END IF;
	--KOTAK DI BAWAH M
		IF B_BAWAH >= G27_ATAS AND B_BAWAH <= G27_BAWAH AND B_KIRI < G27_KANAN AND B_KANAN > G27_KIRI THEN
			B_ATAS := G27_ATAS - 30;
			B_BAWAH := G27_ATAS;
			END IF;
	--GARIS HORIZONTAL_3 DI BAWAH M
		IF B_BAWAH >= G31_ATAS AND B_BAWAH <= G31_BAWAH AND B_KIRI < G31_KANAN AND B_KANAN > G31_KIRI THEN
			B_ATAS := G31_ATAS - 30;
			B_BAWAH := G31_ATAS;
			END IF;
	--GARIS HORIZONTAL DI BAWAH A
		IF B_BAWAH >= G32_ATAS AND B_BAWAH <= G32_BAWAH AND B_KIRI < G32_KANAN AND B_KANAN > G32_KIRI THEN
			B_ATAS := G32_ATAS - 30;
			B_BAWAH := G32_ATAS;
			END IF;
	--KOTAK DI BAWAH A
		IF B_BAWAH >= G33_ATAS AND B_BAWAH <= G33_BAWAH AND B_KIRI < G33_KANAN AND B_KANAN > G33_KIRI THEN
			B_ATAS := G33_ATAS - 30;
			B_BAWAH := G33_ATAS;
			END IF;
	--GARIS HORIZONTAL_1 DI BAWAH U
		IF B_BAWAH >= G42_ATAS AND B_BAWAH <= G42_BAWAH AND B_KIRI < G42_KANAN AND B_KANAN > G42_KIRI THEN
			B_ATAS := G42_ATAS - 30;
			B_BAWAH := G42_ATAS;
			END IF;
	--GARIS HORIZONTAL_3 DI BAWAH U
		IF B_BAWAH >= G44_ATAS AND B_BAWAH <= G44_BAWAH AND B_KIRI < G44_KANAN AND B_KANAN > G44_KIRI THEN
			B_ATAS := G44_ATAS - 30;
			B_BAWAH := G44_ATAS;
			END IF;
	--GARIS HORIZONTAL_4 DI BAWAH U
		IF B_BAWAH >= G45_ATAS AND B_BAWAH <= G45_BAWAH AND B_KIRI < G45_KANAN AND B_KANAN > G45_KIRI THEN
			B_ATAS := G45_ATAS - 30;
			B_BAWAH := G45_ATAS;
			END IF;
	--GARIS HORIZONTAL_5 DI BAWAH U
		IF B_BAWAH >= G46_ATAS AND B_BAWAH <= G46_BAWAH AND B_KIRI < G46_KANAN AND B_KANAN > G46_KIRI THEN
			B_ATAS := G46_ATAS - 30;
			B_BAWAH := G46_ATAS;
			END IF;
	--TELEPORT 1
		IF B_KANAN <= G47_KANAN AND B_KIRI >= G47_KIRI AND B_ATAS >= G47_ATAS AND B_BAWAH <= G47_BAWAH THEN
			B_ATAS := 130;
			B_BAWAH := 130 + 30;
			B_KIRI := 160;
			B_KANAN := 160 + 30;
			END IF;
	--TELEPORT 2
		IF B_KANAN <= G48_KANAN AND B_KIRI >= G48_KIRI AND B_ATAS >= G48_ATAS AND B_BAWAH <= G48_BAWAH THEN
			B_ATAS := 10;
			B_BAWAH := 10 + 30;
			B_KIRI := 10;
			B_KANAN := 10 + 30;
			END IF;
	--TELEPORT 4
		IF B_KANAN <= G50_KANAN AND B_KIRI >= G50_KIRI AND B_ATAS >= G50_ATAS AND B_BAWAH <= G50_BAWAH THEN
			B_ATAS := 170;
			B_BAWAH := 170 + 30;
			B_KIRI := 10;
			B_KANAN := 10 + 30;
			END IF;
	--TELEPORT 5
		IF B_KANAN <= G51_KANAN AND B_KIRI >= G51_KIRI AND B_ATAS >= G51_ATAS AND B_BAWAH <= G51_BAWAH THEN
			B_ATAS := 230;
			B_BAWAH := 230 + 30;
			B_KIRI := 320;
			B_KANAN := 320 + 30;
			END IF;
	--TELEPORT 6
		IF B_KANAN <= G52_KANAN AND B_KIRI >= G52_KIRI AND B_ATAS >= G52_ATAS AND B_BAWAH <= G52_BAWAH THEN
			B_ATAS := 170;
			B_BAWAH := 170 + 30;
			B_KIRI := 320;
			B_KANAN := 320 + 30;
			END IF;
			
	ELSIF clock40hz'event and clock40hz = '1' AND i_M_US = '1' AND i_K_US = '1' AND i_H_US = '0' AND i_M_BT = '1' THEN
		B_KANAN		:= B_KANAN + KECEPATAN;  ---Arah kanan
		B_KIRI 		:= B_KIRI + KECEPATAN;
		
		IF B_KANAN >= 639 THEN
			B_KANAN := 639;
			B_KIRI := 639 -49;
			END IF;
			
	--BINGKAI KANAN
		IF B_KANAN >= G4_KIRI THEN
			B_KANAN := G4_KIRI;
			B_KIRI := G4_KIRI - 30;
			END IF;
	--GARIS VERTIKAL ANTARA I DAN M
		IF B_KANAN >= G5_KIRI AND B_KANAN <= G5_KANAN AND B_ATAS < G5_BAWAH THEN
			B_KANAN := G5_KIRI;
			B_KIRI := G5_KIRI - 30;
			END IF;
	--GARIS VERTIKAL M_1
		IF B_KANAN >= G7_KIRI AND B_KANAN <= G7_KANAN AND B_BAWAH > G7_ATAS AND B_ATAS < G7_BAWAH THEN
			B_KANAN := G7_KIRI;
			B_KIRI := G7_KIRI - 30;
			END IF;
	--GARIS VERTIKAL M_2 AMPE BAWAH
		IF B_KANAN >= G8_KIRI AND B_KANAN <= G8_KANAN AND B_BAWAH > G8_ATAS THEN
			B_KANAN := G8_KIRI;
			B_KIRI := G8_KIRI - 30;
			END IF;
	--GARIS VERTIKAL M_3
		IF B_KANAN >= G9_KIRI AND B_KANAN <= G9_KANAN AND B_BAWAH > G9_ATAS AND B_ATAS < G9_BAWAH THEN
			B_KANAN := G9_KIRI;
			B_KIRI := G9_KIRI - 30;
			END IF;
	--GARIS VERTIKAL M_4
		IF B_KANAN >= G10_KIRI AND B_KANAN <= G10_KANAN AND B_BAWAH > G10_ATAS AND B_ATAS < G10_BAWAH THEN
			B_KANAN := G10_KIRI;
			B_KIRI := G10_KIRI - 30;
			END IF;
	--GARIS VERTIKAL ANTARA M DAN A
		IF B_KANAN >= G15_KIRI AND B_KANAN <= G15_KANAN AND B_ATAS < G15_BAWAH THEN
			B_KANAN := G15_KIRI;
			B_KIRI := G15_KIRI - 30;
			END IF;
	--KOTAK DI TENGAH A
		IF B_KANAN >= G16_KIRI AND B_KANAN <= G16_KANAN AND B_BAWAH > G16_ATAS AND B_ATAS < G16_BAWAH THEN
			B_KANAN := G16_KIRI;
			B_KIRI := G16_KIRI - 30;
			END IF;
	--KOTAK DI KANAN A
		IF B_KANAN >= G19_KIRI AND B_KANAN <= G19_KANAN AND B_ATAS < G19_BAWAH THEN
			B_KANAN := G19_KIRI;
			B_KIRI := G19_KIRI - 30;
			END IF;
	--GARIS VERTIKAL A_1 AMPE UJUNG BAWAH
		IF B_KANAN >= G20_KIRI AND B_KANAN <= G20_KANAN AND B_BAWAH > G20_ATAS THEN
			B_KANAN := G20_KIRI;
			B_KIRI := G20_KIRI - 30;
			END IF;
	--GARIS VERTIKAL A_2 AMPE LEKUKAN BAWAH
		IF B_KANAN >= G21_KIRI AND B_KANAN <= G21_KANAN AND B_BAWAH > G21_ATAS AND B_ATAS < G21_BAWAH THEN
			B_KANAN := G21_KIRI;
			B_KIRI := G21_KIRI - 30;
			END IF;
	--KOTAK DI BAWAH I
		IF B_KANAN >= G22_KIRI AND B_KANAN <= G22_KANAN AND B_BAWAH > G22_ATAS AND B_ATAS < G22_BAWAH THEN
			B_KANAN := G22_KIRI;
			B_KIRI := G22_KIRI - 30;
			END IF;
	--GARIS HORIZONTAL_1 DI BAWAH M
		IF B_KANAN >= G26_KIRI AND B_KANAN <= G26_KANAN AND B_BAWAH > G26_ATAS AND B_ATAS < G26_BAWAH THEN
			B_KANAN := G26_KIRI;
			B_KIRI := G26_KIRI - 30;
			END IF;
	--GARIS VERTIKAL_1 DI BAWAH M
		IF B_KANAN >= G28_KIRI AND B_KANAN <= G28_KANAN AND B_BAWAH > G28_ATAS AND B_ATAS < G28_BAWAH THEN
			B_KANAN := G28_KIRI;
			B_KIRI := G28_KIRI - 30;
			END IF;
	--GARIS HORIZONTAL_3 DI BAWAH M
		IF B_KANAN >= G31_KIRI AND B_KANAN <= G31_KANAN AND B_BAWAH > G31_ATAS AND B_ATAS < G31_BAWAH THEN
			B_KANAN := G31_KIRI;
			B_KIRI := G31_KIRI - 30;
			END IF;
	--KOTAK DI BAWAH A
		IF B_KANAN >= G33_KIRI AND B_KANAN <= G33_KANAN AND B_BAWAH > G33_ATAS AND B_ATAS < G33_BAWAH THEN
			B_KANAN := G33_KIRI;
			B_KIRI := G33_KIRI - 30;
			END IF;
	--GARIS VERTIKAL DI BAWAH A
		IF B_KANAN >= G34_KIRI AND B_KANAN <= G34_KANAN AND B_BAWAH > G34_ATAS THEN
			B_KANAN := G34_KIRI;
			B_KIRI := G34_KIRI - 30;
			END IF;
	--GARIS VERTIKAL_1 DI KANAN A
		IF B_KANAN >= G35_KIRI AND B_KANAN <= G35_KANAN AND B_ATAS < G35_BAWAH THEN
			B_KANAN := G35_KIRI;
			B_KIRI := G35_KIRI - 30;
			END IF;
	--GARIS VERTIKAL_2 DI KANAN A
		IF B_KANAN >= G36_KIRI AND B_KANAN <= G36_KANAN AND B_ATAS < G36_BAWAH THEN
			B_KANAN := G36_KIRI;
			B_KIRI := G36_KIRI - 30;
			END IF;
	--GARIS VERTIKAL_1 DI BAWAH U
		IF B_KANAN >= G40_KIRI AND B_KANAN <= G40_KANAN AND B_BAWAH > G40_ATAS AND B_ATAS < G40_BAWAH THEN
			B_KANAN := G40_KIRI;
			B_KIRI := G40_KIRI - 30;
			END IF;
	--GARIS VERTIKAL_2 DI BAWAH U
		IF B_KANAN >= G41_KIRI AND B_KANAN <= G41_KANAN AND B_BAWAH > G41_ATAS AND B_ATAS < G41_BAWAH THEN
			B_KANAN := G41_KIRI;
			B_KIRI := G41_KIRI - 30;
			END IF;
	--GARIS HORIZONTAL_4 DI BAWAH U
		IF B_KANAN >= G45_KIRI AND B_KANAN <= G45_KANAN AND B_BAWAH > G45_ATAS AND B_ATAS < G45_BAWAH THEN
			B_KANAN := G45_KIRI;
			B_KIRI := G45_KIRI - 30;
			END IF;
	--TELEPORT 10
		IF B_KANAN <= G56_KANAN AND B_KIRI >= G56_KIRI AND B_ATAS >= G56_ATAS AND B_BAWAH <= G56_BAWAH THEN
			B_ATAS := 130;
			B_BAWAH := 130 + 30;
			B_KIRI := 360;
			B_KANAN := 360 + 30;
			END IF;
	--TELEPORT 13
		IF B_KANAN <= G59_KANAN AND B_KIRI >= G59_KIRI AND B_ATAS >= G59_ATAS AND B_BAWAH <= G59_BAWAH THEN
			B_ATAS := 150;
			B_BAWAH := 150 + 30;
			B_KIRI := 590;
			B_KANAN := 590 + 30;
			END IF;
	
	ELSIF clock40hz'event and clock40hz = '1' AND i_M_US = '1' AND i_K_US = '1' AND i_H_US = '1' AND i_M_BT = '0' THEN
		B_KANAN 	:= B_KANAN - KECEPATAN;  ---Arah Kiri
		B_KIRI 		:= B_KIRI - KECEPATAN;
		
		IF B_KIRI <= 0 THEN
			B_KIRI := 0;
			B_KANAN := 49;
			END IF;
			
	--BINGKAI KIRI
		IF B_KIRI <= G2_KANAN THEN
			B_KIRI := G2_KANAN;
			B_KANAN := G2_KANAN + 30;
			END IF;
	--GARIS VERTIKAL ANTARA I DAN M
		IF B_KIRI <= G5_KANAN AND B_KIRI >= G5_KIRI AND B_ATAS < G5_BAWAH THEN
			B_KIRI := G5_KANAN;
			B_KANAN := G5_KANAN + 30;
			END IF;	
	--GARIS VERTIKAL M_1
		IF B_KIRI <= G7_KANAN AND B_KIRI >= G7_KIRI AND B_ATAS < G7_BAWAH AND B_BAWAH > G7_ATAS THEN
			B_KIRI := G7_KANAN;
			B_KANAN := G7_KANAN + 30;
			END IF;	
	--GARIS VERTIKAL M_2 AMPE BAWAH
		IF B_KIRI <= G8_KANAN AND B_KIRI >= G8_KIRI AND B_BAWAH > G8_ATAS THEN
			B_KIRI := G8_KANAN;
			B_KANAN := G8_KANAN + 30;
			END IF;	
	--GARIS VERTIKAL M_3
		IF B_KIRI <= G9_KANAN AND B_KIRI >= G9_KIRI AND B_ATAS < G9_BAWAH AND B_BAWAH > G9_ATAS THEN
			B_KIRI := G9_KANAN;
			B_KANAN := G9_KANAN + 30;
			END IF;		
	--GARIS VERTIKAL M_4
		IF B_KIRI <= G10_KANAN AND B_KIRI >= G10_KIRI AND B_ATAS < G10_BAWAH AND B_BAWAH > G10_ATAS THEN
			B_KIRI := G10_KANAN;
			B_KANAN := G10_KANAN + 30;
			END IF;		
	--GARIS VERTIKAL ANTARA M DAN A
		IF B_KIRI <= G15_KANAN AND B_KIRI >= G15_KIRI AND B_ATAS < G15_BAWAH THEN
			B_KIRI := G15_KANAN;
			B_KANAN := G15_KANAN + 30;
			END IF;	
	--KOTAK DI TENGAH A
		IF B_KIRI <= G16_KANAN AND B_KIRI >= G16_KIRI AND B_ATAS < G16_BAWAH AND B_BAWAH > G16_ATAS THEN
			B_KIRI := G16_KANAN;
			B_KANAN := G16_KANAN + 30;
			END IF;	
	--KOTAK DI KANAN A
		IF B_KIRI <= G19_KANAN AND B_KIRI >= G19_KIRI AND B_ATAS < G19_BAWAH THEN
			B_KIRI := G19_KANAN;
			B_KANAN := G19_KANAN + 30;
			END IF;	
	--GARIS VERTIKAL A_1 AMPE UJUNG BAWAH
		IF B_KIRI <= G20_KANAN AND B_KIRI >= G20_KIRI AND B_BAWAH > G20_ATAS THEN
			B_KIRI := G20_KANAN;
			B_KANAN := G20_KANAN + 30;
			END IF;	
	--GARIS VERTIKAL A_2 AMPE LEKUKAN BAWAH
		IF B_KIRI <= G21_KANAN AND B_KIRI >= G21_KIRI AND B_ATAS < G21_BAWAH AND B_BAWAH > G21_ATAS THEN
			B_KIRI := G21_KANAN;
			B_KANAN := G21_KANAN + 30;
			END IF;	
	--KOTAK DI BAWAH I
		IF B_KIRI <= G22_KANAN AND B_KIRI >= G22_KIRI AND B_ATAS < G22_BAWAH AND B_BAWAH > G22_ATAS THEN
			B_KIRI := G22_KANAN;
			B_KANAN := G22_KANAN + 30;
			END IF;	
	--GARIS HORIZONTAL_1 DI BAWAH I
		IF B_KIRI <= G23_KANAN AND B_KIRI >= G23_KIRI AND B_ATAS < G23_BAWAH AND B_BAWAH > G23_ATAS THEN
			B_KIRI := G23_KANAN;
			B_KANAN := G23_KANAN + 30;
			END IF;	
	--GARIS HORIZONTAL_3 DI BAWAH I
		IF B_KIRI <= G25_KANAN AND B_KIRI >= G25_KIRI AND B_ATAS < G25_BAWAH AND B_BAWAH > G25_ATAS THEN
			B_KIRI := G25_KANAN;
			B_KANAN := G25_KANAN + 30;
			END IF;	
	--GARIS VERTIKAL_2 DI BAWAH M
		IF B_KIRI <= G29_KANAN AND B_KIRI >= G29_KIRI AND B_ATAS < G29_BAWAH AND B_BAWAH > G29_ATAS THEN
			B_KIRI := G29_KANAN;
			B_KANAN := G29_KANAN + 30;
			END IF;	
	--GARIS HORIZONTAL_2 DI BAWAH M
		IF B_KIRI <= G30_KANAN AND B_KIRI >= G30_KIRI AND B_ATAS < G30_BAWAH AND B_BAWAH > G30_ATAS THEN
			B_KIRI := G30_KANAN;
			B_KANAN := G30_KANAN + 30;
			END IF;
	--GARIS HORIZONTAL DI BAWAH A
		IF B_KIRI <= G32_KANAN AND B_KIRI >= G32_KIRI AND B_ATAS < G32_BAWAH AND B_BAWAH > G32_ATAS THEN
			B_KIRI := G32_KANAN;
			B_KANAN := G32_KANAN + 30;
			END IF;	
	--GARIS VERTIKAL DI BAWAH A
		IF B_KIRI <= G34_KANAN AND B_KIRI >= G34_KIRI AND B_BAWAH > G34_ATAS THEN
			B_KIRI := G34_KANAN;
			B_KANAN := G34_KANAN + 30;
			END IF;	
	--GARIS VERTIKAL_2 DI KANAN A
		IF B_KIRI <= G36_KANAN AND B_KIRI >= G36_KIRI AND B_ATAS < G36_BAWAH AND B_BAWAH > G36_ATAS THEN
			B_KIRI := G36_KANAN;
			B_KANAN := G36_KANAN + 30;
			END IF;
	--GARIS VERTIKAL_1 DI BAWAH U
		IF B_KIRI <= G40_KANAN AND B_KIRI >= G40_KIRI AND B_ATAS < G40_BAWAH AND B_BAWAH > G40_ATAS THEN
			B_KIRI := G40_KANAN;
			B_KANAN := G40_KANAN + 30;
			END IF;	
	--GARIS VERTIKAL_2 DI BAWAH U
		IF B_KIRI <= G41_KANAN AND B_KIRI >= G41_KIRI AND B_ATAS < G41_BAWAH AND B_BAWAH > G41_ATAS THEN
			B_KIRI := G41_KANAN;
			B_KANAN := G41_KANAN + 30;
			END IF;	
	--GARIS HORIZONTAL_3 DI BAWAH U
		IF B_KIRI <= G44_KANAN AND B_KIRI >= G44_KIRI AND B_ATAS < G44_BAWAH AND B_BAWAH > G44_ATAS THEN
			B_KIRI := G44_KANAN;
			B_KANAN := G44_KANAN + 30;
			END IF;	
	--GARIS HORIZONTAL_5 DI BAWAH U
		IF B_KIRI <= G46_KANAN AND B_KIRI >= G46_KIRI AND B_ATAS < G46_BAWAH AND B_BAWAH > G46_ATAS THEN
			B_KIRI := G46_KANAN;
			B_KANAN := G46_KANAN + 30;
			END IF;	
	--TELEPORT 7
		IF B_KANAN <= G53_KANAN AND B_KIRI >= G53_KIRI AND B_ATAS >= G53_ATAS AND B_BAWAH <= G53_BAWAH THEN
			B_ATAS := 10;
			B_BAWAH := 10 + 30;
			B_KIRI := 10;
			B_KANAN := 10 + 30;
			END IF;
	--TELEPORT 8
		IF B_KANAN <= G54_KANAN AND B_KIRI >= G54_KIRI AND B_ATAS >= G54_ATAS AND B_BAWAH <= G54_BAWAH THEN
			B_ATAS := 10;
			B_BAWAH := 10 + 30;
			B_KIRI := 375;
			B_KANAN := 375 + 30;
			END IF;

ELSE

B_KIRI := B_KIRI;
B_KANAN := B_KANAN;
B_BAWAH := B_BAWAH;
B_ATAS := B_ATAS;

END IF;

	--WARNA PEMBATAS LEVEL 2
	IF ((i_pixel_column > B_KIRI) AND (i_pixel_column < B_KANAN) AND (i_pixel_row >B_ATAS) AND (i_pixel_row < B_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"00"; o_blue <= X"00";
			
		ELSIF ((i_pixel_column > G1_KIRI) AND (i_pixel_column < G1_KANAN) AND (i_pixel_row > G1_ATAS) AND (i_pixel_row < G1_BAWAH)) THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G2_KIRI) AND (i_pixel_column < G2_KANAN) AND (i_pixel_row > G2_ATAS) AND (i_pixel_row < G2_BAWAH)) THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G3_KIRI) AND (i_pixel_column < G3_KANAN) AND (i_pixel_row > G3_ATAS) AND (i_pixel_row < G3_BAWAH)) THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G4_KIRI) AND (i_pixel_column < G4_KANAN) AND (i_pixel_row > G4_ATAS) AND (i_pixel_row < G4_BAWAH)) THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G5_KIRI) AND (i_pixel_column < G5_KANAN) AND (i_pixel_row > G5_ATAS) AND (i_pixel_row < G5_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G6_KIRI) AND (i_pixel_column < G6_KANAN) AND (i_pixel_row > G6_ATAS) AND (i_pixel_row < G6_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G7_KIRI) AND (i_pixel_column < G7_KANAN) AND (i_pixel_row > G7_ATAS) AND (i_pixel_row < G7_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G8_KIRI) AND (i_pixel_column < G8_KANAN) AND (i_pixel_row > G8_ATAS) AND (i_pixel_row < G8_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";
		ELSIF ((i_pixel_column > G9_KIRI) AND (i_pixel_column < G9_KANAN) AND (i_pixel_row > G9_ATAS) AND (i_pixel_row < G9_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G10_KIRI) AND (i_pixel_column < G10_KANAN) AND (i_pixel_row > G10_ATAS) AND (i_pixel_row < G10_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G11_KIRI) AND (i_pixel_column < G11_KANAN) AND (i_pixel_row > G11_ATAS) AND (i_pixel_row < G11_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G12_KIRI) AND (i_pixel_column < G12_KANAN) AND (i_pixel_row > G12_ATAS) AND (i_pixel_row < G12_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G13_KIRI) AND (i_pixel_column < G13_KANAN) AND (i_pixel_row > G13_ATAS) AND (i_pixel_row < G13_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G14_KIRI) AND (i_pixel_column < G14_KANAN) AND (i_pixel_row > G14_ATAS) AND (i_pixel_row < G14_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G15_KIRI) AND (i_pixel_column < G15_KANAN) AND (i_pixel_row > G15_ATAS) AND (i_pixel_row < G15_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G16_KIRI) AND (i_pixel_column < G16_KANAN) AND (i_pixel_row > G16_ATAS) AND (i_pixel_row < G16_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G17_KIRI) AND (i_pixel_column < G17_KANAN) AND (i_pixel_row > G17_ATAS) AND (i_pixel_row < G17_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G18_KIRI) AND (i_pixel_column < G18_KANAN) AND (i_pixel_row > G18_ATAS) AND (i_pixel_row < G18_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G19_KIRI) AND (i_pixel_column < G19_KANAN) AND (i_pixel_row > G19_ATAS) AND (i_pixel_row < G19_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G20_KIRI) AND (i_pixel_column < G20_KANAN) AND (i_pixel_row > G20_ATAS) AND (i_pixel_row < G20_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G21_KIRI) AND (i_pixel_column < G21_KANAN) AND (i_pixel_row > G21_ATAS) AND (i_pixel_row < G21_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G22_KIRI) AND (i_pixel_column < G22_KANAN) AND (i_pixel_row > G22_ATAS) AND (i_pixel_row < G22_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G23_KIRI) AND (i_pixel_column < G23_KANAN) AND (i_pixel_row > G23_ATAS) AND (i_pixel_row < G23_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G24_KIRI) AND (i_pixel_column < G24_KANAN) AND (i_pixel_row > G24_ATAS) AND (i_pixel_row < G24_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G25_KIRI) AND (i_pixel_column < G25_KANAN) AND (i_pixel_row > G25_ATAS) AND (i_pixel_row < G25_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G26_KIRI) AND (i_pixel_column < G26_KANAN) AND (i_pixel_row > G26_ATAS) AND (i_pixel_row < G26_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G27_KIRI) AND (i_pixel_column < G27_KANAN) AND (i_pixel_row > G27_ATAS) AND (i_pixel_row < G27_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G28_KIRI) AND (i_pixel_column < G28_KANAN) AND (i_pixel_row > G28_ATAS) AND (i_pixel_row < G28_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G29_KIRI) AND (i_pixel_column < G29_KANAN) AND (i_pixel_row > G29_ATAS) AND (i_pixel_row < G29_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G30_KIRI) AND (i_pixel_column < G30_KANAN) AND (i_pixel_row > G30_ATAS) AND (i_pixel_row < G30_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G31_KIRI) AND (i_pixel_column < G31_KANAN) AND (i_pixel_row > G31_ATAS) AND (i_pixel_row < G31_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G32_KIRI) AND (i_pixel_column < G32_KANAN) AND (i_pixel_row > G32_ATAS) AND (i_pixel_row < G32_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G33_KIRI) AND (i_pixel_column < G33_KANAN) AND (i_pixel_row > G33_ATAS) AND (i_pixel_row < G33_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G34_KIRI) AND (i_pixel_column < G34_KANAN) AND (i_pixel_row > G34_ATAS) AND (i_pixel_row < G34_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G35_KIRI) AND (i_pixel_column < G35_KANAN) AND (i_pixel_row > G35_ATAS) AND (i_pixel_row < G35_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G36_KIRI) AND (i_pixel_column < G36_KANAN) AND (i_pixel_row > G36_ATAS) AND (i_pixel_row < G36_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G37_KIRI) AND (i_pixel_column < G37_KANAN) AND (i_pixel_row > G37_ATAS) AND (i_pixel_row < G37_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G40_KIRI) AND (i_pixel_column < G40_KANAN) AND (i_pixel_row > G40_ATAS) AND (i_pixel_row < G40_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G41_KIRI) AND (i_pixel_column < G41_KANAN) AND (i_pixel_row > G41_ATAS) AND (i_pixel_row < G41_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G42_KIRI) AND (i_pixel_column < G42_KANAN) AND (i_pixel_row > G42_ATAS) AND (i_pixel_row < G42_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";		
		ELSIF ((i_pixel_column > G44_KIRI) AND (i_pixel_column < G44_KANAN) AND (i_pixel_row > G44_ATAS) AND (i_pixel_row < G44_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G45_KIRI) AND (i_pixel_column < G45_KANAN) AND (i_pixel_row > G45_ATAS) AND (i_pixel_row < G45_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G46_KIRI) AND (i_pixel_column < G46_KANAN) AND (i_pixel_row > G46_ATAS) AND (i_pixel_row < G46_BAWAH)) AND B_ATAS >= P_ATAS AND B_KIRI >= P_KIRI AND B_KANAN <= P_KANAN AND B_BAWAH <= P_BAWAH THEN
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";	
		ELSIF ((i_pixel_column > G47_KIRI) AND (i_pixel_column < G47_KANAN) AND (i_pixel_row > G47_ATAS) AND (i_pixel_row < G47_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G48_KIRI) AND (i_pixel_column < G48_KANAN) AND (i_pixel_row > G48_ATAS) AND (i_pixel_row < G48_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G49_KIRI) AND (i_pixel_column < G49_KANAN) AND (i_pixel_row > G49_ATAS) AND (i_pixel_row < G49_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G50_KIRI) AND (i_pixel_column < G50_KANAN) AND (i_pixel_row > G50_ATAS) AND (i_pixel_row < G50_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";		
		ELSIF ((i_pixel_column > G51_KIRI) AND (i_pixel_column < G51_KANAN) AND (i_pixel_row > G51_ATAS) AND (i_pixel_row < G51_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G52_KIRI) AND (i_pixel_column < G52_KANAN) AND (i_pixel_row > G52_ATAS) AND (i_pixel_row < G52_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G53_KIRI) AND (i_pixel_column < G53_KANAN) AND (i_pixel_row > G53_ATAS) AND (i_pixel_row < G53_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G54_KIRI) AND (i_pixel_column < G54_KANAN) AND (i_pixel_row > G54_ATAS) AND (i_pixel_row < G54_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G55_KIRI) AND (i_pixel_column < G55_KANAN) AND (i_pixel_row > G55_ATAS) AND (i_pixel_row < G55_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G56_KIRI) AND (i_pixel_column < G56_KANAN) AND (i_pixel_row > G56_ATAS) AND (i_pixel_row < G56_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G57_KIRI) AND (i_pixel_column < G57_KANAN) AND (i_pixel_row > G57_ATAS) AND (i_pixel_row < G57_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G58_KIRI) AND (i_pixel_column < G58_KANAN) AND (i_pixel_row > G58_ATAS) AND (i_pixel_row < G58_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G59_KIRI) AND (i_pixel_column < G59_KANAN) AND (i_pixel_row > G59_ATAS) AND (i_pixel_row < G59_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G60_KIRI) AND (i_pixel_column < G60_KANAN) AND (i_pixel_row > G60_ATAS) AND (i_pixel_row < G60_BAWAH)) THEN
			o_red <= X"C8"; o_green <= X"C8"; o_blue <= X"C8";	
		ELSIF ((i_pixel_column > G61_KIRI) AND (i_pixel_column < G61_KANAN) AND (i_pixel_row > G61_ATAS) AND (i_pixel_row < G61_BAWAH)) THEN
			o_red <= X"64"; o_green <= X"FA"; o_blue <= X"C8";
	
	--PERUBAHAN WARNA PEMBATAS LEVEL 2
		ELSIF ((i_pixel_column > G5_KIRI) AND (i_pixel_column < G5_KANAN) AND (i_pixel_row > G5_ATAS) AND (i_pixel_row < G5_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G6_KIRI) AND (i_pixel_column < G6_KANAN) AND (i_pixel_row > G6_ATAS) AND (i_pixel_row < G6_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G7_KIRI) AND (i_pixel_column < G7_KANAN) AND (i_pixel_row > G7_ATAS) AND (i_pixel_row < G7_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G8_KIRI) AND (i_pixel_column < G8_KANAN) AND (i_pixel_row > G8_ATAS) AND (i_pixel_row < G8_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G9_KIRI) AND (i_pixel_column < G9_KANAN) AND (i_pixel_row > G9_ATAS) AND (i_pixel_row < G9_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G10_KIRI) AND (i_pixel_column < G10_KANAN) AND (i_pixel_row > G10_ATAS) AND (i_pixel_row < G10_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G11_KIRI) AND (i_pixel_column < G11_KANAN) AND (i_pixel_row > G11_ATAS) AND (i_pixel_row < G11_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G12_KIRI) AND (i_pixel_column < G12_KANAN) AND (i_pixel_row > G12_ATAS) AND (i_pixel_row < G12_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G13_KIRI) AND (i_pixel_column < G13_KANAN) AND (i_pixel_row > G13_ATAS) AND (i_pixel_row < G13_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G14_KIRI) AND (i_pixel_column < G14_KANAN) AND (i_pixel_row > G14_ATAS) AND (i_pixel_row < G14_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G15_KIRI) AND (i_pixel_column < G15_KANAN) AND (i_pixel_row > G15_ATAS) AND (i_pixel_row < G15_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G16_KIRI) AND (i_pixel_column < G16_KANAN) AND (i_pixel_row > G16_ATAS) AND (i_pixel_row < G16_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G17_KIRI) AND (i_pixel_column < G17_KANAN) AND (i_pixel_row > G17_ATAS) AND (i_pixel_row < G17_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G18_KIRI) AND (i_pixel_column < G18_KANAN) AND (i_pixel_row > G18_ATAS) AND (i_pixel_row < G18_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G19_KIRI) AND (i_pixel_column < G19_KANAN) AND (i_pixel_row > G19_ATAS) AND (i_pixel_row < G19_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G20_KIRI) AND (i_pixel_column < G20_KANAN) AND (i_pixel_row > G20_ATAS) AND (i_pixel_row < G20_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G21_KIRI) AND (i_pixel_column < G21_KANAN) AND (i_pixel_row > G21_ATAS) AND (i_pixel_row < G21_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G22_KIRI) AND (i_pixel_column < G22_KANAN) AND (i_pixel_row > G22_ATAS) AND (i_pixel_row < G22_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G23_KIRI) AND (i_pixel_column < G23_KANAN) AND (i_pixel_row > G23_ATAS) AND (i_pixel_row < G23_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G24_KIRI) AND (i_pixel_column < G24_KANAN) AND (i_pixel_row > G24_ATAS) AND (i_pixel_row < G24_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G25_KIRI) AND (i_pixel_column < G25_KANAN) AND (i_pixel_row > G25_ATAS) AND (i_pixel_row < G25_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G26_KIRI) AND (i_pixel_column < G26_KANAN) AND (i_pixel_row > G26_ATAS) AND (i_pixel_row < G26_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G27_KIRI) AND (i_pixel_column < G27_KANAN) AND (i_pixel_row > G27_ATAS) AND (i_pixel_row < G27_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G28_KIRI) AND (i_pixel_column < G28_KANAN) AND (i_pixel_row > G28_ATAS) AND (i_pixel_row < G28_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G29_KIRI) AND (i_pixel_column < G29_KANAN) AND (i_pixel_row > G29_ATAS) AND (i_pixel_row < G29_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G30_KIRI) AND (i_pixel_column < G30_KANAN) AND (i_pixel_row > G30_ATAS) AND (i_pixel_row < G30_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G31_KIRI) AND (i_pixel_column < G31_KANAN) AND (i_pixel_row >G31_ATAS) AND (i_pixel_row < G31_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G32_KIRI) AND (i_pixel_column < G32_KANAN) AND (i_pixel_row > G32_ATAS) AND (i_pixel_row < G32_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G33_KIRI) AND (i_pixel_column < G33_KANAN) AND (i_pixel_row > G33_ATAS) AND (i_pixel_row < G33_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G34_KIRI) AND (i_pixel_column < G34_KANAN) AND (i_pixel_row > G34_ATAS) AND (i_pixel_row < G34_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G35_KIRI) AND (i_pixel_column < G35_KANAN) AND (i_pixel_row > G35_ATAS) AND (i_pixel_row < G35_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G36_KIRI) AND (i_pixel_column < G36_KANAN) AND (i_pixel_row > G36_ATAS) AND (i_pixel_row < G36_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G37_KIRI) AND (i_pixel_column < G37_KANAN) AND (i_pixel_row > G37_ATAS) AND (i_pixel_row < G37_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G40_KIRI) AND (i_pixel_column < G40_KANAN) AND (i_pixel_row > G40_ATAS) AND (i_pixel_row < G40_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G41_KIRI) AND (i_pixel_column < G41_KANAN) AND (i_pixel_row > G41_ATAS) AND (i_pixel_row < G41_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G42_KIRI) AND (i_pixel_column < G42_KANAN) AND (i_pixel_row > G42_ATAS) AND (i_pixel_row < G42_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G44_KIRI) AND (i_pixel_column < G44_KANAN) AND (i_pixel_row > G44_ATAS) AND (i_pixel_row < G44_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G45_KIRI) AND (i_pixel_column < G45_KANAN) AND (i_pixel_row > G45_ATAS) AND (i_pixel_row < G45_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G46_KIRI) AND (i_pixel_column < G46_KANAN) AND (i_pixel_row > G46_ATAS) AND (i_pixel_row < G46_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		
		--WAKTU
		ELSIF ((i_pixel_column > G63_KIRI) AND (i_pixel_column < G63_KANAN) AND (i_pixel_row > G63_ATAS) AND (i_pixel_row < G63_BAWAH)) THEN
			o_red <= X"00"; o_green <= X"FF"; o_blue <= X"00";
		ELSIF ((i_pixel_column > G63A_KIRI) AND (i_pixel_column < G63A_KANAN) AND (i_pixel_row > G63A_ATAS) AND (i_pixel_row < G63A_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"00";
		ELSIF ((i_pixel_column > G63B_KIRI) AND (i_pixel_column < G63B_KANAN) AND (i_pixel_row > G63B_ATAS) AND (i_pixel_row < G63B_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"00"; o_blue <= X"00";
		ELSE 
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
	END IF;
END IF;

--MENANG KALAH
IF i_K_BT = '1' AND MENANG = TRUE THEN --TAMPILAN MENANG
	IF ((i_pixel_column > G120_KIRI) AND (i_pixel_column < G120_KANAN) AND (i_pixel_row > G120_ATAS) AND (i_pixel_row < G120_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G121_KIRI) AND (i_pixel_column < G121_KANAN) AND (i_pixel_row > G121_ATAS) AND (i_pixel_row < G121_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G122_KIRI) AND (i_pixel_column < G122_KANAN) AND (i_pixel_row > G122_ATAS) AND (i_pixel_row < G122_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G123_KIRI) AND (i_pixel_column < G123_KANAN) AND (i_pixel_row > G123_ATAS) AND (i_pixel_row < G123_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G124_KIRI) AND (i_pixel_column < G124_KANAN) AND (i_pixel_row > G124_ATAS) AND (i_pixel_row < G124_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";		
		ELSIF ((i_pixel_column > G125_KIRI) AND (i_pixel_column < G125_KANAN) AND (i_pixel_row > G125_ATAS) AND (i_pixel_row < G125_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G126_KIRI) AND (i_pixel_column < G126_KANAN) AND (i_pixel_row > G126_ATAS) AND (i_pixel_row < G126_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G127_KIRI) AND (i_pixel_column < G127_KANAN) AND (i_pixel_row > G127_ATAS) AND (i_pixel_row < G127_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G128_KIRI) AND (i_pixel_column < G128_KANAN) AND (i_pixel_row > G128_ATAS) AND (i_pixel_row < G128_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G129_KIRI) AND (i_pixel_column < G129_KANAN) AND (i_pixel_row > G129_ATAS) AND (i_pixel_row < G129_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G130_KIRI) AND (i_pixel_column < G130_KANAN) AND (i_pixel_row > G130_ATAS) AND (i_pixel_row < G130_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G131_KIRI) AND (i_pixel_column < G131_KANAN) AND (i_pixel_row > G131_ATAS) AND (i_pixel_row < G131_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		
		ELSE
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";
	END IF;
	
ELSIF i_K_BT = '1' AND (KALAH = TRUE OR KALAH1 = TRUE) THEN --TAMPILAN KALAH
	IF ((i_pixel_column > G105_KIRI) AND (i_pixel_column < G105_KANAN) AND (i_pixel_row > G105_ATAS) AND (i_pixel_row < G105_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G106_KIRI) AND (i_pixel_column < G106_KANAN) AND (i_pixel_row > G106_ATAS) AND (i_pixel_row < G106_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G107_KIRI) AND (i_pixel_column < G107_KANAN) AND (i_pixel_row > G107_ATAS) AND (i_pixel_row < G107_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G108_KIRI) AND (i_pixel_column < G108_KANAN) AND (i_pixel_row > G108_ATAS) AND (i_pixel_row < G108_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";		
		ELSIF ((i_pixel_column > G109_KIRI) AND (i_pixel_column < G109_KANAN) AND (i_pixel_row > G109_ATAS) AND (i_pixel_row < G109_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G110_KIRI) AND (i_pixel_column < G110_KANAN) AND (i_pixel_row > G110_ATAS) AND (i_pixel_row < G110_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G111_KIRI) AND (i_pixel_column < G111_KANAN) AND (i_pixel_row > G111_ATAS) AND (i_pixel_row < G111_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G112_KIRI) AND (i_pixel_column < G112_KANAN) AND (i_pixel_row > G112_ATAS) AND (i_pixel_row < G112_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G113_KIRI) AND (i_pixel_column < G113_KANAN) AND (i_pixel_row > G113_ATAS) AND (i_pixel_row < G113_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G114_KIRI) AND (i_pixel_column < G114_KANAN) AND (i_pixel_row > G114_ATAS) AND (i_pixel_row < G114_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G115_KIRI) AND (i_pixel_column < G115_KANAN) AND (i_pixel_row > G115_ATAS) AND (i_pixel_row < G115_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G116_KIRI) AND (i_pixel_column < G116_KANAN) AND (i_pixel_row > G116_ATAS) AND (i_pixel_row < G116_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
		ELSIF ((i_pixel_column > G117_KIRI) AND (i_pixel_column < G117_KANAN) AND (i_pixel_row > G117_ATAS) AND (i_pixel_row < G117_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G118_KIRI) AND (i_pixel_column < G118_KANAN) AND (i_pixel_row > G118_ATAS) AND (i_pixel_row < G118_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";	
		ELSIF ((i_pixel_column > G119_KIRI) AND (i_pixel_column < G119_KANAN) AND (i_pixel_row > G119_ATAS) AND (i_pixel_row < G119_BAWAH)) THEN
			o_red <= X"FF"; o_green <= X"FF"; o_blue <= X"FF";
			
		ELSE
			o_red <= X"00"; o_green <= X"00"; o_blue <= X"00";
		END IF;
	END IF;

--RESTART
IF RESTART = TRUE THEN
	MENANG		:= FALSE;
	KALAH		:= FALSE;
	KALAH1		:= FALSE;
	G63_ATAS	:= 10;
	G63A_ATAS	:= 10;
	G63B_ATAS	:= 10;
	B_ATAS		:= 10; 
	B_KIRI 		:= 20; 
	B_KANAN 	:= 50; 
	B_BAWAH		:= 40;
	G62_ATAS	:= 10;
	G62A_ATAS	:= 10;
	G62B_ATAS	:= 10;
	B1_ATAS		:= 10; 
	B1_KIRI		:= 10; 
	B1_KANAN 	:= 60; 
	B1_BAWAH 	:= 60;
END IF;

--PENGAKTIFAN RESTART
IF i_K_BT = '0' AND i_M_US = '0' THEN
	RESTART	:= TRUE;
	ELSE
		RESTART	:= FALSE;
END IF;

--RESET
IF RESET = TRUE THEN
	LEVEL		:= 1;
	MENANG		:= FALSE;
	KALAH		:= FALSE;
	KALAH1		:= FALSE;
	G63_ATAS	:= 10;
	G63A_ATAS	:= 10;
	G63B_ATAS	:= 10;
	B_ATAS		:= 10; 
	B_KIRI 		:= 20; 
	B_KANAN 	:= 50; 
	B_BAWAH		:= 40;
	G62_ATAS	:= 10;
	G62A_ATAS	:= 10;
	G62B_ATAS	:= 10;
	B1_ATAS		:= 10; 
	B1_KIRI		:= 10; 
	B1_KANAN 	:= 60; 
	B1_BAWAH 	:= 60;
END IF;

--PENGAKTIFAN RESET
IF i_K_BT = '0' AND i_K_US = '0' THEN
	RESET	:= TRUE;
	ELSE
		RESET := FALSE;
END IF;

END PROCESS;

tempik : clockdiv
	PORT MAP ( 
				CLK => i_H_BT,
				DIVOUT => clock40hz
			);

END behavioral; 